module log2_32b ( a, result);
  input  [31:0] a ;
  output wire [31:0] result ;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
    n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
    n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
    n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
    n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
    n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
    n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
    n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
    n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
    n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
    n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
    n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
    n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
    n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
    n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
    n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
    n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
    n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
    n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
    n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
    n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
    n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
    n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
    n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
    n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
    n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
    n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
    n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
    n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
    n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
    n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
    n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
    n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
    n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
    n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
    n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
    n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
    n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
    n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
    n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
    n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
    n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
    n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
    n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
    n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
    n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
    n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
    n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
    n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
    n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
    n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
    n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
    n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
    n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
    n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
    n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
    n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
    n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
    n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
    n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
    n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
    n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
    n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
    n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
    n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
    n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
    n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
    n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
    n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
    n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
    n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
    n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
    n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
    n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
    n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
    n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
    n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
    n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
    n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
    n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
    n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
    n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
    n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
    n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
    n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
    n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
    n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
    n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
    n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
    n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
    n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
    n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
    n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
    n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
    n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
    n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
    n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
    n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
    n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
    n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
    n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
    n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
    n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
    n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
    n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
    n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
    n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
    n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
    n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
    n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
    n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
    n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
    n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
    n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
    n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
    n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
    n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
    n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
    n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
    n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
    n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
    n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
    n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
    n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
    n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
    n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
    n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
    n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
    n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
    n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
    n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
    n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
    n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
    n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
    n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
    n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
    n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
    n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
    n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
    n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
    n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
    n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
    n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
    n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
    n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
    n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
    n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
    n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
    n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
    n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
    n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
    n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
    n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
    n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
    n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
    n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
    n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
    n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
    n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
    n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
    n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
    n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
    n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
    n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
    n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
    n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
    n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
    n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
    n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
    n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
    n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
    n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
    n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
    n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
    n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
    n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
    n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
    n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
    n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
    n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
    n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
    n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
    n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
    n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
    n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
    n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
    n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
    n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
    n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
    n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
    n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
    n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
    n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
    n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
    n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
    n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
    n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
    n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
    n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
    n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
    n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
    n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
    n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
    n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
    n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
    n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
    n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
    n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
    n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
    n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
    n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
    n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
    n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
    n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
    n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
    n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
    n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
    n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
    n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
    n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
    n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
    n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
    n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
    n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
    n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
    n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
    n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
    n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
    n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
    n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
    n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
    n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
    n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
    n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
    n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
    n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
    n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
    n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
    n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
    n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
    n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
    n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
    n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
    n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
    n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
    n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
    n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
    n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
    n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
    n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
    n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
    n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
    n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
    n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
    n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
    n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
    n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
    n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
    n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
    n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
    n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
    n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
    n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
    n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
    n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
    n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
    n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
    n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
    n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
    n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
    n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
    n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
    n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
    n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
    n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
    n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
    n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
    n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
    n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
    n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
    n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
    n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
    n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
    n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
    n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
    n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
    n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
    n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
    n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
    n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
    n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
    n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
    n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
    n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
    n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
    n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
    n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
    n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
    n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
    n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
    n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
    n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
    n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
    n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
    n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
    n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
    n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
    n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
    n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
    n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
    n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
    n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
    n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
    n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
    n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
    n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
    n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
    n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
    n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
    n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
    n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
    n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
    n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
    n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
    n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
    n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
    n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
    n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
    n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
    n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
    n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
    n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
    n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
    n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
    n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
    n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
    n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
    n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
    n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
    n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
    n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
    n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
    n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
    n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
    n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
    n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
    n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
    n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
    n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
    n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
    n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
    n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
    n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
    n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
    n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
    n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
    n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
    n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
    n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
    n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
    n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
    n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
    n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
    n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
    n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
    n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
    n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
    n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
    n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
    n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
    n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
    n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
    n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
    n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
    n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
    n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
    n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
    n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
    n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
    n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
    n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
    n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
    n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
    n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
    n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
    n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
    n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
    n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
    n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
    n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
    n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
    n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
    n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
    n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
    n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
    n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
    n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
    n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
    n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
    n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
    n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
    n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
    n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
    n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
    n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
    n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
    n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
    n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
    n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
    n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
    n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
    n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
    n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
    n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
    n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
    n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
    n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
    n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
    n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
    n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
    n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
    n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
    n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
    n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
    n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
    n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
    n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
    n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
    n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
    n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
    n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
    n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
    n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
    n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
    n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
    n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
    n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
    n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
    n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
    n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
    n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
    n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
    n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
    n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
    n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
    n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
    n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
    n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
    n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
    n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
    n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
    n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
    n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
    n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
    n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
    n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
    n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
    n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
    n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
    n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
    n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
    n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
    n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
    n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
    n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
    n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
    n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
    n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
    n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
    n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
    n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
    n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
    n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
    n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
    n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
    n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
    n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
    n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
    n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
    n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
    n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
    n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
    n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
    n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
    n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
    n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
    n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
    n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
    n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
    n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
    n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
    n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
    n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
    n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
    n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
    n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
    n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
    n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
    n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
    n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
    n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
    n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
    n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
    n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
    n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
    n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
    n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
    n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
    n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
    n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
    n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
    n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
    n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
    n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
    n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
    n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
    n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
    n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
    n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
    n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
    n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
    n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
    n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
    n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
    n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
    n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
    n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
    n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
    n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
    n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
    n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
    n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
    n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
    n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
    n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
    n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
    n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
    n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
    n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
    n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
    n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
    n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
    n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
    n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
    n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
    n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
    n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
    n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
    n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
    n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
    n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
    n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
    n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
    n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
    n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
    n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
    n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
    n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
    n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
    n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
    n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
    n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
    n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
    n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
    n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
    n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
    n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
    n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
    n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
    n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
    n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
    n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
    n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
    n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
    n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
    n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
    n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
    n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
    n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
    n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
    n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
    n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
    n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
    n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
    n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
    n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
    n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
    n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
    n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
    n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
    n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
    n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
    n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
    n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
    n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
    n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
    n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
    n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
    n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
    n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
    n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
    n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
    n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
    n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
    n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
    n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
    n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
    n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
    n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
    n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
    n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
    n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
    n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
    n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
    n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
    n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
    n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
    n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
    n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
    n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
    n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
    n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
    n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
    n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
    n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
    n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
    n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
    n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
    n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
    n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
    n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
    n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
    n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
    n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
    n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
    n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
    n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
    n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
    n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
    n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
    n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
    n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
    n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
    n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
    n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
    n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
    n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
    n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
    n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
    n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
    n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
    n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
    n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
    n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
    n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
    n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
    n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
    n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
    n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
    n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
    n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
    n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
    n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
    n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
    n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
    n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
    n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
    n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
    n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
    n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
    n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
    n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
    n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
    n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
    n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
    n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
    n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
    n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
    n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
    n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
    n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
    n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
    n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
    n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
    n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
    n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
    n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
    n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
    n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
    n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
    n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
    n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
    n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
    n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
    n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
    n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
    n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
    n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
    n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
    n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
    n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
    n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
    n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
    n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
    n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
    n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
    n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
    n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
    n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
    n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
    n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
    n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
    n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
    n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
    n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
    n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
    n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
    n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
    n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
    n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
    n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
    n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
    n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
    n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
    n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
    n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
    n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
    n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
    n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
    n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
    n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
    n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
    n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
    n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
    n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
    n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
    n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
    n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
    n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
    n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
    n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
    n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
    n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
    n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
    n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
    n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
    n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
    n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
    n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
    n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
    n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
    n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
    n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
    n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
    n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
    n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
    n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
    n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
    n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
    n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
    n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
    n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
    n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
    n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
    n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
    n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
    n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
    n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
    n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
    n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
    n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
    n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
    n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
    n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
    n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
    n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
    n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
    n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
    n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
    n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
    n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
    n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
    n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
    n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
    n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
    n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
    n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
    n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
    n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
    n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
    n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
    n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
    n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
    n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
    n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
    n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
    n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
    n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
    n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
    n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
    n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
    n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
    n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
    n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
    n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
    n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
    n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
    n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
    n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
    n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
    n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
    n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
    n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
    n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
    n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
    n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
    n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
    n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
    n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
    n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
    n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
    n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
    n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
    n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
    n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
    n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
    n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
    n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
    n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
    n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
    n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
    n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
    n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
    n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
    n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
    n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
    n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
    n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
    n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
    n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
    n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
    n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
    n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
    n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
    n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
    n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
    n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
    n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
    n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
    n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
    n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
    n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
    n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
    n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
    n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
    n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
    n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
    n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
    n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
    n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
    n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
    n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
    n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
    n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
    n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
    n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
    n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
    n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
    n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
    n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
    n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
    n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
    n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
    n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
    n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
    n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
    n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
    n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
    n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
    n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
    n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
    n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
    n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
    n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
    n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
    n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
    n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
    n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
    n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
    n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
    n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
    n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
    n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
    n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
    n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
    n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
    n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
    n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
    n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
    n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
    n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
    n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
    n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
    n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
    n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
    n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
    n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
    n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
    n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
    n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
    n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
    n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
    n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
    n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
    n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
    n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
    n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
    n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
    n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
    n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
    n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
    n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
    n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
    n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
    n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
    n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
    n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
    n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
    n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
    n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
    n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
    n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
    n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
    n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
    n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
    n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
    n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
    n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
    n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
    n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
    n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
    n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
    n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
    n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
    n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
    n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
    n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
    n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
    n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
    n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
    n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
    n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
    n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
    n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
    n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
    n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
    n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
    n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
    n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
    n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
    n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
    n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
    n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
    n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
    n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
    n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
    n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
    n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
    n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
    n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
    n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
    n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
    n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
    n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
    n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
    n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
    n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
    n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
    n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
    n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
    n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
    n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
    n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
    n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
    n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
    n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
    n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
    n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
    n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
    n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
    n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
    n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
    n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
    n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
    n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
    n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
    n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
    n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
    n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
    n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
    n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
    n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
    n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
    n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
    n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
    n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
    n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
    n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
    n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
    n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
    n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
    n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
    n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
    n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
    n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
    n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
    n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
    n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
    n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
    n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
    n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
    n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
    n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
    n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
    n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
    n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
    n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
    n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
    n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
    n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
    n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
    n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
    n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
    n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
    n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
    n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
    n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
    n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
    n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
    n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
    n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
    n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
    n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
    n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
    n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
    n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
    n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
    n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
    n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
    n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
    n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
    n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
    n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
    n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
    n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
    n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
    n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
    n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
    n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
    n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
    n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
    n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
    n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
    n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
    n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
    n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
    n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
    n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
    n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
    n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
    n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
    n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
    n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
    n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
    n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
    n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
    n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
    n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
    n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
    n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
    n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
    n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
    n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
    n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
    n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
    n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
    n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
    n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
    n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
    n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
    n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
    n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
    n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
    n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
    n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
    n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
    n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
    n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
    n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
    n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
    n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
    n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
    n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
    n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
    n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
    n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
    n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
    n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
    n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
    n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
    n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
    n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
    n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
    n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
    n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
    n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
    n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
    n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
    n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
    n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
    n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
    n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
    n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
    n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
    n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
    n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
    n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
    n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
    n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
    n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
    n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
    n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
    n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
    n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
    n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
    n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
    n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
    n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
    n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
    n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
    n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
    n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
    n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
    n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
    n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
    n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
    n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
    n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
    n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
    n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
    n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
    n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
    n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
    n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
    n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
    n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
    n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
    n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
    n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
    n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
    n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
    n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
    n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
    n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
    n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
    n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
    n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
    n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
    n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
    n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
    n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324,
    n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
    n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
    n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
    n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
    n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
    n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
    n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
    n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396,
    n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405,
    n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
    n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
    n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
    n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
    n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
    n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
    n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468,
    n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477,
    n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486,
    n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
    n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
    n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
    n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
    n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
    n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540,
    n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549,
    n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558,
    n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
    n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
    n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
    n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612,
    n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630,
    n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
    n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
    n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684,
    n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
    n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
    n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
    n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756,
    n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774,
    n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
    n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
    n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
    n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
    n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828,
    n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837,
    n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846,
    n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
    n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
    n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
    n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
    n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900,
    n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909,
    n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918,
    n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
    n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
    n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
    n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
    n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
    n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972,
    n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
    n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990,
    n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
    n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
    n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
    n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
    n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
    n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044,
    n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053,
    n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
    n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
    n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
    n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
    n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
    n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
    n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116,
    n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
    n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134,
    n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
    n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
    n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
    n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
    n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188,
    n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
    n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
    n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
    n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260,
    n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278,
    n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
    n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
    n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332,
    n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350,
    n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
    n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
    n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
    n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
    n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
    n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404,
    n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
    n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422,
    n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
    n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
    n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
    n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
    n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
    n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476,
    n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
    n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
    n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
    n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
    n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
    n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
    n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
    n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548,
    n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
    n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
    n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
    n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
    n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
    n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
    n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
    n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620,
    n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
    n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
    n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
    n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
    n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
    n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
    n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
    n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692,
    n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
    n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
    n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
    n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,
    n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
    n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
    n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
    n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764,
    n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
    n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782,
    n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
    n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,
    n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
    n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
    n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
    n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836,
    n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
    n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854,
    n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
    n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
    n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
    n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
    n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
    n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908,
    n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
    n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926,
    n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
    n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
    n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
    n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
    n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124,
    n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
    n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
    n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
    n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
    n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
    n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
    n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
    n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
    n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
    n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
    n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268,
    n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
    n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
    n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
    n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
    n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340,
    n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
    n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
    n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
    n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
    n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
    n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
    n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
    n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412,
    n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
    n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430,
    n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
    n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
    n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
    n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
    n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
    n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484,
    n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
    n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
    n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
    n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
    n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
    n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
    n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556,
    n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
    n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
    n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
    n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
    n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
    n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
    n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
    n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628,
    n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
    n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646,
    n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
    n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
    n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
    n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
    n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
    n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700,
    n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
    n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718,
    n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
    n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
    n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
    n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
    n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
    n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772,
    n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
    n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790,
    n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
    n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
    n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
    n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
    n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
    n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844,
    n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853,
    n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862,
    n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
    n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
    n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
    n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
    n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
    n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916,
    n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925,
    n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934,
    n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
    n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
    n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
    n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
    n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
    n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988,
    n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997,
    n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006,
    n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
    n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
    n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
    n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
    n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
    n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060,
    n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069,
    n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078,
    n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
    n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
    n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132,
    n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150,
    n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
    n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
    n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
    n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
    n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204,
    n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
    n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222,
    n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
    n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
    n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
    n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
    n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
    n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276,
    n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
    n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294,
    n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303,
    n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
    n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
    n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
    n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
    n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348,
    n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
    n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366,
    n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
    n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
    n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
    n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
    n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420,
    n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438,
    n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
    n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
    n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
    n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
    n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
    n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
    n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
    n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
    n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
    n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
    n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
    n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654,
    n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
    n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
    n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
    n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
    n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708,
    n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726,
    n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
    n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
    n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
    n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
    n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780,
    n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789,
    n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798,
    n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
    n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
    n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
    n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
    n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
    n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852,
    n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
    n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870,
    n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879,
    n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
    n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
    n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
    n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
    n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924,
    n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933,
    n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942,
    n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
    n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
    n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
    n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
    n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
    n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996,
    n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
    n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
    n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
    n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
    n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
    n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068,
    n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
    n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086,
    n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
    n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
    n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
    n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
    n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140,
    n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158,
    n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
    n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
    n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
    n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
    n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
    n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212,
    n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
    n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230,
    n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
    n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
    n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
    n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
    n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
    n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284,
    n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
    n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302,
    n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
    n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
    n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
    n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
    n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356,
    n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365,
    n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374,
    n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
    n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
    n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
    n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
    n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
    n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428,
    n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437,
    n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446,
    n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
    n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
    n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
    n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
    n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
    n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500,
    n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
    n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518,
    n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
    n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
    n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
    n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
    n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
    n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572,
    n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
    n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590,
    n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
    n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
    n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
    n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
    n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
    n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644,
    n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
    n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662,
    n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
    n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
    n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
    n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
    n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
    n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716,
    n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
    n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734,
    n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
    n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
    n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
    n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
    n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
    n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
    n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878,
    n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
    n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
    n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
    n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
    n26915, n26916, n26917, n26918, n26919, n26920, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
    n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
    n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
    n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
    n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
    n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014,
    n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
    n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
    n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
    n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
    n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
    n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
    n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
    n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
    n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
    n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
    n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
    n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
    n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
    n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
    n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158,
    n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
    n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
    n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
    n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
    n27195, n27196, n27197, n27198, n27200, n27201, n27202, n27203, n27204,
    n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
    n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222,
    n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231,
    n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240,
    n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
    n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
    n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
    n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276,
    n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285,
    n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294,
    n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
    n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
    n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
    n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
    n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
    n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348,
    n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357,
    n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366,
    n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
    n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384,
    n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
    n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
    n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
    n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420,
    n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429,
    n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438,
    n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447,
    n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,
    n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
    n27466, n27467, n27468, n27470, n27471, n27472, n27473, n27474, n27475,
    n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484,
    n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493,
    n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502,
    n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511,
    n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
    n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
    n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
    n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
    n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556,
    n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
    n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574,
    n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
    n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
    n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
    n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
    n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628,
    n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
    n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646,
    n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655,
    n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
    n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
    n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
    n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
    n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700,
    n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
    n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718,
    n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27728,
    n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
    n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
    n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
    n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764,
    n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773,
    n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782,
    n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
    n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800,
    n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
    n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
    n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
    n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836,
    n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845,
    n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854,
    n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
    n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872,
    n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
    n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
    n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
    n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908,
    n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
    n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926,
    n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935,
    n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944,
    n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
    n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
    n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
    n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980,
    n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989,
    n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999,
    n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008,
    n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
    n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
    n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
    n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
    n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053,
    n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062,
    n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071,
    n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080,
    n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
    n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
    n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
    n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
    n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
    n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134,
    n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143,
    n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152,
    n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
    n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
    n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
    n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
    n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
    n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206,
    n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215,
    n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224,
    n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
    n28234, n28235, n28236, n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252,
    n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270,
    n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
    n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
    n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324,
    n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342,
    n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
    n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
    n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
    n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
    n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396,
    n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405,
    n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414,
    n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423,
    n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432,
    n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
    n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
    n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
    n28460, n28461, n28462, n28463, n28464, n28465, n28467, n28468, n28469,
    n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478,
    n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487,
    n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496,
    n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
    n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
    n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
    n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532,
    n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541,
    n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550,
    n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559,
    n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568,
    n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
    n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
    n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
    n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604,
    n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613,
    n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622,
    n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631,
    n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640,
    n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
    n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
    n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
    n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676,
    n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28685, n28686,
    n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695,
    n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704,
    n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
    n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
    n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
    n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740,
    n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749,
    n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758,
    n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767,
    n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776,
    n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
    n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794,
    n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
    n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812,
    n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821,
    n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830,
    n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839,
    n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848,
    n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
    n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866,
    n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
    n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884,
    n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893,
    n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902,
    n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912,
    n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
    n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
    n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
    n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948,
    n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957,
    n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966,
    n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
    n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
    n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
    n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
    n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
    n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020,
    n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029,
    n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038,
    n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047,
    n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056,
    n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
    n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
    n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
    n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092,
    n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101,
    n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110,
    n29111, n29112, n29113, n29115, n29116, n29117, n29118, n29119, n29120,
    n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
    n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
    n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
    n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156,
    n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165,
    n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
    n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
    n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192,
    n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
    n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
    n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
    n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228,
    n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237,
    n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
    n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
    n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
    n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
    n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
    n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
    n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300,
    n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309,
    n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29318, n29319,
    n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328,
    n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
    n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346,
    n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
    n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364,
    n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373,
    n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382,
    n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391,
    n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400,
    n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
    n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
    n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
    n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436,
    n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445,
    n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454,
    n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463,
    n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472,
    n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
    n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490,
    n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
    n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508,
    n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517,
    n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526,
    n29527, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
    n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
    n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554,
    n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
    n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572,
    n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581,
    n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590,
    n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599,
    n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608,
    n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
    n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
    n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
    n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644,
    n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653,
    n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
    n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671,
    n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
    n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
    n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
    n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
    n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716,
    n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725,
    n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
    n29735, n29736, n29737, n29738, n29739, n29741, n29742, n29743, n29744,
    n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
    n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
    n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
    n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780,
    n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789,
    n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
    n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807,
    n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
    n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
    n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
    n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
    n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852,
    n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861,
    n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
    n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879,
    n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
    n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
    n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
    n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
    n29916, n29917, n29918, n29919, n29920, n29921, n29923, n29924, n29925,
    n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934,
    n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943,
    n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952,
    n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
    n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970,
    n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
    n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988,
    n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997,
    n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006,
    n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015,
    n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
    n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
    n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
    n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
    n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060,
    n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069,
    n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
    n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087,
    n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096,
    n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
    n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
    n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
    n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
    n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
    n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
    n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196,
    n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205,
    n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
    n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
    n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
    n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
    n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
    n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
    n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268,
    n30269, n30270, n30271, n30272, n30274, n30275, n30276, n30277, n30278,
    n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287,
    n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296,
    n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
    n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314,
    n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
    n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332,
    n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341,
    n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350,
    n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359,
    n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368,
    n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
    n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386,
    n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
    n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404,
    n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413,
    n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
    n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431,
    n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30441,
    n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450,
    n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
    n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468,
    n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477,
    n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
    n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495,
    n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
    n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
    n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522,
    n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
    n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540,
    n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549,
    n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
    n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567,
    n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576,
    n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
    n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594,
    n30595, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604,
    n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613,
    n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
    n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
    n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
    n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
    n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658,
    n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
    n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676,
    n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685,
    n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694,
    n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
    n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712,
    n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
    n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730,
    n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
    n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748,
    n30749, n30750, n30751, n30753, n30754, n30755, n30756, n30757, n30758,
    n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
    n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
    n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
    n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
    n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
    n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812,
    n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821,
    n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
    n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839,
    n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848,
    n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
    n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866,
    n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
    n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884,
    n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893,
    n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903,
    n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912,
    n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
    n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930,
    n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
    n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948,
    n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957,
    n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966,
    n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975,
    n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984,
    n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
    n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002,
    n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
    n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020,
    n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029,
    n31030, n31031, n31033, n31034, n31035, n31036, n31037, n31038, n31039,
    n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048,
    n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
    n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066,
    n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
    n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084,
    n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093,
    n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102,
    n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
    n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
    n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
    n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138,
    n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
    n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156,
    n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165,
    n31166, n31167, n31168, n31169, n31171, n31172, n31173, n31174, n31175,
    n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
    n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
    n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202,
    n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
    n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220,
    n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229,
    n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238,
    n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
    n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
    n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
    n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274,
    n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
    n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
    n31293, n31294, n31296, n31297, n31298, n31299, n31300, n31301, n31302,
    n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311,
    n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320,
    n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
    n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
    n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
    n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356,
    n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365,
    n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374,
    n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383,
    n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392,
    n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
    n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410,
    n31411, n31412, n31413, n31415, n31416, n31417, n31418, n31419, n31420,
    n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429,
    n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438,
    n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
    n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
    n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
    n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474,
    n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
    n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492,
    n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501,
    n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510,
    n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
    n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31529,
    n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538,
    n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
    n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556,
    n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565,
    n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574,
    n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583,
    n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
    n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
    n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
    n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
    n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628,
    n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31638,
    n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647,
    n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656,
    n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
    n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674,
    n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683,
    n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692,
    n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701,
    n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710,
    n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
    n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728,
    n31729, n31730, n31731, n31732, n31733, n31734, n31736, n31737, n31738,
    n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
    n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
    n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765,
    n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774,
    n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
    n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792,
    n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
    n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810,
    n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819,
    n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828,
    n31829, n31830, n31831, n31832, n31834, n31835, n31836, n31837, n31838,
    n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
    n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856,
    n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
    n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874,
    n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883,
    n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892,
    n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901,
    n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910,
    n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
    n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
    n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938,
    n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
    n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956,
    n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965,
    n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974,
    n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
    n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992,
    n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32002,
    n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
    n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
    n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029,
    n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038,
    n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047,
    n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056,
    n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
    n32066, n32067, n32068, n32069, n32070, n32072, n32073, n32074, n32075,
    n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084,
    n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093,
    n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102,
    n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111,
    n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
    n32121, n32122, n32123;
  assign n65 =  a[4]  & ~ a[5] ;
  assign n66 = ~ a[4]  &  a[5] ;
  assign n67 = ~n65 & ~n66;
  assign n68 =  a[2]  & ~ a[3] ;
  assign n69 = ~ a[2]  &  a[3] ;
  assign n70 = ~n68 & ~n69;
  assign n71 = n67 & ~n70;
  assign n72 = ~ a[29]  &  a[30] ;
  assign n73 =  a[29]  & ~ a[30] ;
  assign n74 = ~n72 & ~n73;
  assign n75 =  a[31]  & ~n74;
  assign n76 = ~ a[24]  & ~ a[25] ;
  assign n77 = ~ a[23]  &  a[26] ;
  assign n78 = n76 & n77;
  assign n79 =  a[27]  &  a[28] ;
  assign n80 = n73 & n79;
  assign n81 = n78 & n80;
  assign n82 = ~ a[27]  & ~ a[28] ;
  assign n83 = n73 & n82;
  assign n84 =  a[24]  &  a[25] ;
  assign n85 = n77 & n84;
  assign n86 = n83 & n85;
  assign n87 = ~ a[23]  & ~ a[26] ;
  assign n88 = n76 & n87;
  assign n89 =  a[29]  &  a[30] ;
  assign n90 = n79 & n89;
  assign n91 = n88 & n90;
  assign n92 =  a[23]  & ~ a[26] ;
  assign n93 = ~ a[24]  &  a[25] ;
  assign n94 = n92 & n93;
  assign n95 = n83 & n94;
  assign n96 = n84 & n92;
  assign n97 = ~ a[29]  & ~ a[30] ;
  assign n98 = n82 & n97;
  assign n99 = n96 & n98;
  assign n100 = ~n95 & ~n99;
  assign n101 = n87 & n93;
  assign n102 = n90 & n101;
  assign n103 =  a[27]  & ~ a[28] ;
  assign n104 = n89 & n103;
  assign n105 =  a[23]  &  a[26] ;
  assign n106 = n93 & n105;
  assign n107 = n104 & n106;
  assign n108 = ~n102 & ~n107;
  assign n109 = ~ a[27]  &  a[28] ;
  assign n110 = n72 & n109;
  assign n111 = n96 & n110;
  assign n112 =  a[24]  & ~ a[25] ;
  assign n113 = n92 & n112;
  assign n114 = n72 & n103;
  assign n115 = n113 & n114;
  assign n116 = ~n111 & ~n115;
  assign n117 = n82 & n89;
  assign n118 = n94 & n117;
  assign n119 = n83 & n106;
  assign n120 = ~n118 & ~n119;
  assign n121 = n88 & n117;
  assign n122 = n87 & n112;
  assign n123 = n110 & n122;
  assign n124 = n77 & n93;
  assign n125 = n83 & n124;
  assign n126 = n105 & n112;
  assign n127 = n83 & n126;
  assign n128 = ~n125 & ~n127;
  assign n129 = n97 & n109;
  assign n130 = n113 & n129;
  assign n131 = n76 & n92;
  assign n132 = n129 & n131;
  assign n133 = ~n130 & ~n132;
  assign n134 = n72 & n82;
  assign n135 = n113 & n134;
  assign n136 = n110 & n126;
  assign n137 = ~n135 & ~n136;
  assign n138 = n133 & n137;
  assign n139 = n128 & n138;
  assign n140 = ~n123 & n139;
  assign n141 = ~n121 & n140;
  assign n142 = n98 & n126;
  assign n143 = n79 & n97;
  assign n144 = n122 & n143;
  assign n145 = n78 & n143;
  assign n146 = n104 & n126;
  assign n147 = n78 & n117;
  assign n148 = n77 & n112;
  assign n149 = n117 & n148;
  assign n150 = n114 & n124;
  assign n151 = n114 & n122;
  assign n152 = n101 & n134;
  assign n153 = n72 & n79;
  assign n154 = n126 & n153;
  assign n155 = n117 & n124;
  assign n156 = ~n154 & ~n155;
  assign n157 = n94 & n129;
  assign n158 = n83 & n148;
  assign n159 = ~n157 & ~n158;
  assign n160 = n73 & n109;
  assign n161 = n94 & n160;
  assign n162 = n84 & n105;
  assign n163 = n129 & n162;
  assign n164 = n85 & n143;
  assign n165 = n124 & n143;
  assign n166 = n97 & n103;
  assign n167 = n124 & n166;
  assign n168 = n114 & n126;
  assign n169 = n85 & n153;
  assign n170 = n129 & n148;
  assign n171 = n114 & n131;
  assign n172 = ~n170 & ~n171;
  assign n173 = n88 & n143;
  assign n174 = n89 & n109;
  assign n175 = n106 & n174;
  assign n176 = n84 & n87;
  assign n177 = n117 & n176;
  assign n178 = ~n175 & ~n177;
  assign n179 = ~n173 & n178;
  assign n180 = n172 & n179;
  assign n181 = ~n169 & n180;
  assign n182 = ~n168 & n181;
  assign n183 = ~n167 & n182;
  assign n184 = ~n165 & n183;
  assign n185 = ~n164 & n184;
  assign n186 = ~n163 & n185;
  assign n187 = ~n161 & n186;
  assign n188 = n80 & n124;
  assign n189 = n106 & n114;
  assign n190 = n122 & n153;
  assign n191 = n98 & n162;
  assign n192 = n101 & n166;
  assign n193 = ~n191 & ~n192;
  assign n194 = n110 & n113;
  assign n195 = n193 & ~n194;
  assign n196 = ~n190 & n195;
  assign n197 = ~n189 & n196;
  assign n198 = ~n188 & n197;
  assign n199 = n73 & n103;
  assign n200 = n176 & n199;
  assign n201 = n126 & n199;
  assign n202 = ~n200 & ~n201;
  assign n203 = n126 & n174;
  assign n204 = n202 & ~n203;
  assign n205 = n94 & n143;
  assign n206 = n90 & n148;
  assign n207 = ~n205 & ~n206;
  assign n208 = n204 & n207;
  assign n209 = n198 & n208;
  assign n210 = n187 & n209;
  assign n211 = n159 & n210;
  assign n212 = n156 & n211;
  assign n213 = ~n152 & n212;
  assign n214 = ~n151 & n213;
  assign n215 = ~n150 & n214;
  assign n216 = ~n149 & n215;
  assign n217 = ~n147 & n216;
  assign n218 = ~n146 & n217;
  assign n219 = ~n145 & n218;
  assign n220 = ~n144 & n219;
  assign n221 = ~n142 & n220;
  assign n222 = n80 & n85;
  assign n223 = n117 & n162;
  assign n224 = n85 & n134;
  assign n225 = n88 & n199;
  assign n226 = n94 & n104;
  assign n227 = ~n225 & ~n226;
  assign n228 = n90 & n122;
  assign n229 = n78 & n153;
  assign n230 = ~n228 & ~n229;
  assign n231 = n80 & n106;
  assign n232 = n126 & n134;
  assign n233 = n78 & n174;
  assign n234 = ~n232 & ~n233;
  assign n235 = ~n231 & n234;
  assign n236 = n85 & n110;
  assign n237 = n148 & n199;
  assign n238 = ~n236 & ~n237;
  assign n239 = n85 & n117;
  assign n240 = n143 & n148;
  assign n241 = ~n239 & ~n240;
  assign n242 = n153 & n176;
  assign n243 = n143 & n176;
  assign n244 = ~n242 & ~n243;
  assign n245 = n98 & n124;
  assign n246 = n126 & n166;
  assign n247 = ~n245 & ~n246;
  assign n248 = n104 & n162;
  assign n249 = n80 & n131;
  assign n250 = ~n248 & ~n249;
  assign n251 = n83 & n131;
  assign n252 = n106 & n199;
  assign n253 = ~n251 & ~n252;
  assign n254 = n114 & n176;
  assign n255 = n106 & n134;
  assign n256 = ~n254 & ~n255;
  assign n257 = n253 & n256;
  assign n258 = n250 & n257;
  assign n259 = n247 & n258;
  assign n260 = n244 & n259;
  assign n261 = n241 & n260;
  assign n262 = n238 & n261;
  assign n263 = n235 & n262;
  assign n264 = n230 & n263;
  assign n265 = n227 & n264;
  assign n266 = ~n224 & n265;
  assign n267 = ~n223 & n266;
  assign n268 = ~n222 & n267;
  assign n269 = n76 & n105;
  assign n270 = n80 & n269;
  assign n271 = n83 & n88;
  assign n272 = n131 & n199;
  assign n273 = n126 & n129;
  assign n274 = n131 & n143;
  assign n275 = n113 & n117;
  assign n276 = n110 & n131;
  assign n277 = n96 & n160;
  assign n278 = n134 & n162;
  assign n279 = ~n277 & ~n278;
  assign n280 = n101 & n114;
  assign n281 = n96 & n134;
  assign n282 = ~n280 & ~n281;
  assign n283 = n98 & n131;
  assign n284 = n134 & n148;
  assign n285 = ~n283 & ~n284;
  assign n286 = n131 & n166;
  assign n287 = n90 & n94;
  assign n288 = ~n286 & ~n287;
  assign n289 = n94 & n134;
  assign n290 = n96 & n104;
  assign n291 = ~n289 & ~n290;
  assign n292 = n104 & n131;
  assign n293 = n83 & n162;
  assign n294 = ~n292 & ~n293;
  assign n295 = n124 & n160;
  assign n296 = n94 & n166;
  assign n297 = ~n295 & ~n296;
  assign n298 = n98 & n176;
  assign n299 = n117 & n131;
  assign n300 = ~n298 & ~n299;
  assign n301 = n110 & n176;
  assign n302 = n90 & n124;
  assign n303 = ~n301 & ~n302;
  assign n304 = n88 & n160;
  assign n305 = n104 & n269;
  assign n306 = n129 & n269;
  assign n307 = ~n305 & ~n306;
  assign n308 = ~n304 & n307;
  assign n309 = n303 & n308;
  assign n310 = n300 & n309;
  assign n311 = n297 & n310;
  assign n312 = n294 & n311;
  assign n313 = n291 & n312;
  assign n314 = n288 & n313;
  assign n315 = n285 & n314;
  assign n316 = n282 & n315;
  assign n317 = n279 & n316;
  assign n318 = ~n276 & n317;
  assign n319 = ~n275 & n318;
  assign n320 = ~n274 & n319;
  assign n321 = ~n273 & n320;
  assign n322 = ~n272 & n321;
  assign n323 = ~n271 & n322;
  assign n324 = ~n270 & n323;
  assign n325 = n83 & n101;
  assign n326 = n90 & n162;
  assign n327 = n162 & n174;
  assign n328 = n88 & n114;
  assign n329 = n78 & n134;
  assign n330 = n94 & n153;
  assign n331 = n162 & n166;
  assign n332 = n160 & n269;
  assign n333 = ~n331 & ~n332;
  assign n334 = n174 & n176;
  assign n335 = n94 & n114;
  assign n336 = ~n334 & ~n335;
  assign n337 = n80 & n101;
  assign n338 = n85 & n199;
  assign n339 = n101 & n174;
  assign n340 = n113 & n160;
  assign n341 = ~n339 & ~n340;
  assign n342 = ~n338 & n341;
  assign n343 = ~n337 & n342;
  assign n344 = n336 & n343;
  assign n345 = n333 & n344;
  assign n346 = ~n330 & n345;
  assign n347 = ~n329 & n346;
  assign n348 = ~n328 & n347;
  assign n349 = ~n327 & n348;
  assign n350 = ~n326 & n349;
  assign n351 = ~n325 & n350;
  assign n352 = n122 & n174;
  assign n353 = n134 & n176;
  assign n354 = n124 & n134;
  assign n355 = n134 & n269;
  assign n356 = ~n354 & ~n355;
  assign n357 = n90 & n269;
  assign n358 = n83 & n269;
  assign n359 = ~n357 & ~n358;
  assign n360 = n356 & n359;
  assign n361 = ~n353 & n360;
  assign n362 = ~n352 & n361;
  assign n363 = n80 & n94;
  assign n364 = n110 & n162;
  assign n365 = ~n363 & ~n364;
  assign n366 = n96 & n199;
  assign n367 = n104 & n113;
  assign n368 = n98 & n113;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~n366 & n369;
  assign n371 = n85 & n160;
  assign n372 = n88 & n98;
  assign n373 = ~n371 & ~n372;
  assign n374 = n90 & n96;
  assign n375 = n78 & n129;
  assign n376 = ~n374 & ~n375;
  assign n377 = n373 & n376;
  assign n378 = n370 & n377;
  assign n379 = n365 & n378;
  assign n380 = n362 & n379;
  assign n381 = n351 & n380;
  assign n382 = n324 & n381;
  assign n383 = n268 & n382;
  assign n384 = n221 & n383;
  assign n385 = n141 & n384;
  assign n386 = n120 & n385;
  assign n387 = n116 & n386;
  assign n388 = n108 & n387;
  assign n389 = n100 & n388;
  assign n390 = ~n91 & n389;
  assign n391 = ~n86 & n390;
  assign n392 = ~n81 & n391;
  assign n393 = n85 & n129;
  assign n394 = n124 & n129;
  assign n395 = n90 & n113;
  assign n396 = n78 & n104;
  assign n397 = n106 & n110;
  assign n398 = n131 & n153;
  assign n399 = ~n327 & ~n398;
  assign n400 = n88 & n104;
  assign n401 = ~n335 & ~n400;
  assign n402 = n101 & n104;
  assign n403 = n104 & n148;
  assign n404 = ~n402 & ~n403;
  assign n405 = ~n375 & n404;
  assign n406 = n401 & n405;
  assign n407 = n399 & n406;
  assign n408 = ~n111 & n407;
  assign n409 = ~n397 & n408;
  assign n410 = ~n177 & n409;
  assign n411 = ~n299 & n410;
  assign n412 = ~n396 & n411;
  assign n413 = ~n395 & n412;
  assign n414 = ~n325 & n413;
  assign n415 = ~n293 & n414;
  assign n416 = n78 & n90;
  assign n417 = n117 & n122;
  assign n418 = ~n364 & ~n417;
  assign n419 = n96 & n117;
  assign n420 = n106 & n153;
  assign n421 = ~n419 & ~n420;
  assign n422 = n98 & n148;
  assign n423 = ~n146 & ~n422;
  assign n424 = n101 & n143;
  assign n425 = n166 & n269;
  assign n426 = n114 & n148;
  assign n427 = n110 & n148;
  assign n428 = n80 & n176;
  assign n429 = n80 & n148;
  assign n430 = n148 & n166;
  assign n431 = ~n144 & ~n430;
  assign n432 = ~n201 & n431;
  assign n433 = ~n429 & n432;
  assign n434 = ~n428 & n433;
  assign n435 = n117 & n269;
  assign n436 = n160 & n176;
  assign n437 = ~n435 & ~n436;
  assign n438 = n88 & n166;
  assign n439 = ~n371 & ~n438;
  assign n440 = n437 & n439;
  assign n441 = n434 & n440;
  assign n442 = ~n427 & n441;
  assign n443 = ~n194 & n442;
  assign n444 = ~n426 & n443;
  assign n445 = ~n280 & n444;
  assign n446 = ~n367 & n445;
  assign n447 = ~n425 & n446;
  assign n448 = ~n424 & n447;
  assign n449 = n80 & n122;
  assign n450 = ~n271 & ~n449;
  assign n451 = n199 & n269;
  assign n452 = n85 & n98;
  assign n453 = n98 & n101;
  assign n454 = ~n452 & ~n453;
  assign n455 = ~n289 & n454;
  assign n456 = ~n292 & n455;
  assign n457 = ~n286 & n456;
  assign n458 = ~n225 & n457;
  assign n459 = ~n451 & n458;
  assign n460 = n104 & n176;
  assign n461 = n85 & n104;
  assign n462 = n148 & n153;
  assign n463 = ~n461 & ~n462;
  assign n464 = ~n460 & n463;
  assign n465 = ~n283 & n464;
  assign n466 = n96 & n143;
  assign n467 = ~n233 & ~n466;
  assign n468 = n106 & n129;
  assign n469 = n94 & n110;
  assign n470 = n94 & n199;
  assign n471 = ~n366 & ~n470;
  assign n472 = ~n469 & n471;
  assign n473 = ~n468 & n472;
  assign n474 = n101 & n160;
  assign n475 = ~n188 & ~n474;
  assign n476 = n473 & n475;
  assign n477 = n467 & n476;
  assign n478 = n465 & n477;
  assign n479 = n459 & n478;
  assign n480 = n450 & n479;
  assign n481 = n448 & n480;
  assign n482 = n159 & n481;
  assign n483 = n423 & n482;
  assign n484 = n421 & n483;
  assign n485 = n418 & n484;
  assign n486 = ~n254 & n485;
  assign n487 = ~n416 & n486;
  assign n488 = ~n337 & n487;
  assign n489 = n83 & n176;
  assign n490 = n90 & n106;
  assign n491 = ~n489 & ~n490;
  assign n492 = n166 & n176;
  assign n493 = n129 & n176;
  assign n494 = ~n167 & ~n493;
  assign n495 = n85 & n174;
  assign n496 = n78 & n166;
  assign n497 = ~n495 & ~n496;
  assign n498 = n494 & n497;
  assign n499 = ~n242 & n498;
  assign n500 = ~n189 & n499;
  assign n501 = ~n290 & n500;
  assign n502 = ~n492 & n501;
  assign n503 = ~n231 & n502;
  assign n504 = n143 & n162;
  assign n505 = n96 & n166;
  assign n506 = n96 & n174;
  assign n507 = ~n81 & ~n506;
  assign n508 = ~n275 & ~n334;
  assign n509 = n101 & n153;
  assign n510 = ~n135 & ~n509;
  assign n511 = n114 & n269;
  assign n512 = ~n248 & ~n511;
  assign n513 = n104 & n124;
  assign n514 = n174 & n269;
  assign n515 = ~n306 & ~n357;
  assign n516 = ~n161 & n515;
  assign n517 = ~n332 & n516;
  assign n518 = n96 & n153;
  assign n519 = n122 & n160;
  assign n520 = ~n518 & ~n519;
  assign n521 = n517 & n520;
  assign n522 = ~n514 & n521;
  assign n523 = ~n513 & n522;
  assign n524 = ~n274 & n523;
  assign n525 = n160 & n162;
  assign n526 = ~n272 & ~n525;
  assign n527 = n104 & n122;
  assign n528 = ~n115 & ~n305;
  assign n529 = ~n527 & n528;
  assign n530 = ~n127 & ~n223;
  assign n531 = n101 & n199;
  assign n532 = n148 & n160;
  assign n533 = ~n340 & ~n532;
  assign n534 = ~n531 & n533;
  assign n535 = ~n338 & n534;
  assign n536 = n78 & n98;
  assign n537 = n98 & n122;
  assign n538 = ~n368 & ~n537;
  assign n539 = ~n536 & n538;
  assign n540 = ~n298 & n539;
  assign n541 = ~n358 & n540;
  assign n542 = n535 & n541;
  assign n543 = n530 & n542;
  assign n544 = n529 & n543;
  assign n545 = n526 & n544;
  assign n546 = n524 & n545;
  assign n547 = n512 & n546;
  assign n548 = n510 & n547;
  assign n549 = n508 & n548;
  assign n550 = n507 & n549;
  assign n551 = n108 & n550;
  assign n552 = ~n169 & n551;
  assign n553 = ~n147 & n552;
  assign n554 = ~n505 & n553;
  assign n555 = ~n504 & n554;
  assign n556 = ~n245 & n555;
  assign n557 = n88 & n134;
  assign n558 = n88 & n110;
  assign n559 = ~n557 & ~n558;
  assign n560 = ~n226 & n559;
  assign n561 = ~n277 & n560;
  assign n562 = n80 & n162;
  assign n563 = n85 & n166;
  assign n564 = n78 & n160;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n562 & n565;
  assign n567 = n98 & n269;
  assign n568 = n122 & n166;
  assign n569 = n83 & n122;
  assign n570 = ~n568 & ~n569;
  assign n571 = n88 & n174;
  assign n572 = n570 & ~n571;
  assign n573 = ~n567 & n572;
  assign n574 = n566 & n573;
  assign n575 = n561 & n574;
  assign n576 = n556 & n575;
  assign n577 = n503 & n576;
  assign n578 = n491 & n577;
  assign n579 = n488 & n578;
  assign n580 = n415 & n579;
  assign n581 = n193 & n580;
  assign n582 = ~n152 & n581;
  assign n583 = ~n302 & n582;
  assign n584 = ~n243 & n583;
  assign n585 = ~n394 & n584;
  assign n586 = ~n393 & n585;
  assign n587 = ~n249 & n586;
  assign n588 = ~n392 & ~n587;
  assign n589 = n96 & n129;
  assign n590 = ~n188 & ~n222;
  assign n591 = ~n194 & ~n490;
  assign n592 = n124 & n199;
  assign n593 = ~n228 & ~n592;
  assign n594 = n117 & n126;
  assign n595 = ~n205 & ~n594;
  assign n596 = n593 & n595;
  assign n597 = ~n136 & n596;
  assign n598 = ~n177 & n597;
  assign n599 = ~n394 & n598;
  assign n600 = ~n119 & n599;
  assign n601 = n106 & n143;
  assign n602 = n114 & n162;
  assign n603 = n101 & n129;
  assign n604 = ~n493 & ~n603;
  assign n605 = n359 & n604;
  assign n606 = ~n602 & n605;
  assign n607 = ~n299 & n606;
  assign n608 = ~n107 & n607;
  assign n609 = ~n243 & n608;
  assign n610 = ~n601 & n609;
  assign n611 = ~n393 & n610;
  assign n612 = ~n470 & n611;
  assign n613 = ~n272 & n612;
  assign n614 = ~n340 & n613;
  assign n615 = ~n151 & ~n327;
  assign n616 = ~n229 & n376;
  assign n617 = n110 & n269;
  assign n618 = ~n171 & ~n617;
  assign n619 = n124 & n174;
  assign n620 = n131 & n134;
  assign n621 = ~n619 & ~n620;
  assign n622 = ~n175 & ~n525;
  assign n623 = n162 & n199;
  assign n624 = ~n135 & ~n152;
  assign n625 = ~n335 & n624;
  assign n626 = ~n150 & n625;
  assign n627 = ~n248 & n626;
  assign n628 = ~n164 & n627;
  assign n629 = ~n623 & n628;
  assign n630 = ~n532 & n629;
  assign n631 = ~n86 & n630;
  assign n632 = ~n102 & ~n242;
  assign n633 = n80 & n126;
  assign n634 = ~n424 & ~n633;
  assign n635 = ~n154 & n634;
  assign n636 = ~n400 & n635;
  assign n637 = n101 & n117;
  assign n638 = ~n571 & ~n637;
  assign n639 = n90 & n126;
  assign n640 = ~n505 & ~n639;
  assign n641 = n78 & n114;
  assign n642 = ~n492 & ~n641;
  assign n643 = n640 & n642;
  assign n644 = n638 & n643;
  assign n645 = n636 & n644;
  assign n646 = n632 & n645;
  assign n647 = n631 & n646;
  assign n648 = n622 & n647;
  assign n649 = n621 & n648;
  assign n650 = n618 & n649;
  assign n651 = ~n398 & n650;
  assign n652 = ~n149 & n651;
  assign n653 = ~n223 & n652;
  assign n654 = ~n123 & ~n125;
  assign n655 = n80 & n113;
  assign n656 = n94 & n174;
  assign n657 = n113 & n199;
  assign n658 = ~n452 & ~n657;
  assign n659 = ~n427 & n658;
  assign n660 = ~n353 & n659;
  assign n661 = ~n426 & n660;
  assign n662 = ~n656 & n661;
  assign n663 = ~n292 & n662;
  assign n664 = ~n655 & n663;
  assign n665 = ~n283 & ~n567;
  assign n666 = n83 & n96;
  assign n667 = n153 & n162;
  assign n668 = ~n281 & ~n667;
  assign n669 = ~n430 & n668;
  assign n670 = ~n519 & n669;
  assign n671 = ~n666 & n670;
  assign n672 = n106 & n160;
  assign n673 = n143 & n269;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n144 & ~n568;
  assign n676 = n674 & n675;
  assign n677 = n671 & n676;
  assign n678 = n665 & n677;
  assign n679 = n664 & n678;
  assign n680 = n654 & n679;
  assign n681 = n450 & n680;
  assign n682 = ~n330 & n681;
  assign n683 = ~n419 & n682;
  assign n684 = ~n461 & n683;
  assign n685 = ~n527 & n684;
  assign n686 = ~n422 & n685;
  assign n687 = ~n170 & n686;
  assign n688 = ~n562 & n687;
  assign n689 = n113 & n143;
  assign n690 = ~n190 & ~n689;
  assign n691 = ~n329 & ~n339;
  assign n692 = ~n420 & ~n536;
  assign n693 = ~n468 & n692;
  assign n694 = ~n145 & ~n254;
  assign n695 = n693 & n694;
  assign n696 = n691 & n695;
  assign n697 = n690 & n696;
  assign n698 = n688 & n697;
  assign n699 = n653 & n698;
  assign n700 = n616 & n699;
  assign n701 = n333 & n700;
  assign n702 = n615 & n701;
  assign n703 = n614 & n702;
  assign n704 = n600 & n703;
  assign n705 = n591 & n704;
  assign n706 = n202 & n705;
  assign n707 = n590 & n706;
  assign n708 = ~n514 & n707;
  assign n709 = ~n326 & n708;
  assign n710 = ~n589 & n709;
  assign n711 = ~n587 & ~n710;
  assign n712 = n78 & n199;
  assign n713 = n122 & n134;
  assign n714 = n126 & n143;
  assign n715 = n90 & n131;
  assign n716 = n113 & n166;
  assign n717 = n137 & ~n462;
  assign n718 = ~n367 & n717;
  assign n719 = ~n716 & n718;
  assign n720 = ~n164 & ~n251;
  assign n721 = ~n155 & ~n469;
  assign n722 = ~n374 & n721;
  assign n723 = ~n147 & ~n460;
  assign n724 = n722 & n723;
  assign n725 = ~n355 & n724;
  assign n726 = ~n146 & n725;
  assign n727 = ~n286 & n726;
  assign n728 = ~n567 & n727;
  assign n729 = ~n393 & n728;
  assign n730 = ~n338 & n729;
  assign n731 = ~n145 & ~n571;
  assign n732 = ~n371 & ~n474;
  assign n733 = ~n173 & ~n519;
  assign n734 = ~n158 & n733;
  assign n735 = ~n536 & ~n656;
  assign n736 = n734 & n735;
  assign n737 = n732 & n736;
  assign n738 = ~n242 & n737;
  assign n739 = ~n289 & n738;
  assign n740 = ~n305 & n739;
  assign n741 = ~n248 & n740;
  assign n742 = ~n453 & n741;
  assign n743 = ~n394 & n742;
  assign n744 = ~n95 & n743;
  assign n745 = ~n363 & n744;
  assign n746 = n101 & n110;
  assign n747 = ~n206 & ~n302;
  assign n748 = ~n746 & n747;
  assign n749 = ~n425 & n748;
  assign n750 = ~n99 & n749;
  assign n751 = ~n592 & n750;
  assign n752 = n124 & n153;
  assign n753 = ~n154 & ~n752;
  assign n754 = ~n563 & n753;
  assign n755 = n193 & ~n490;
  assign n756 = ~n237 & n755;
  assign n757 = ~n304 & n756;
  assign n758 = n754 & n757;
  assign n759 = n751 & n758;
  assign n760 = n745 & n759;
  assign n761 = n731 & n760;
  assign n762 = n730 & n761;
  assign n763 = n720 & n762;
  assign n764 = n719 & n763;
  assign n765 = n227 & n764;
  assign n766 = ~n203 & n765;
  assign n767 = ~n715 & n766;
  assign n768 = ~n714 & n767;
  assign n769 = ~n165 & n768;
  assign n770 = ~n429 & n769;
  assign n771 = n80 & n88;
  assign n772 = ~n451 & ~n771;
  assign n773 = ~n190 & ~n240;
  assign n774 = ~n358 & ~n402;
  assign n775 = ~n364 & ~n427;
  assign n776 = ~n278 & ~n328;
  assign n777 = n85 & n90;
  assign n778 = ~n337 & ~n777;
  assign n779 = n776 & n778;
  assign n780 = n775 & n779;
  assign n781 = n774 & n780;
  assign n782 = n773 & n781;
  assign n783 = ~n290 & n782;
  assign n784 = ~n357 & n783;
  assign n785 = ~n416 & n784;
  assign n786 = ~n372 & n785;
  assign n787 = ~n271 & n786;
  assign n788 = ~n86 & ~n493;
  assign n789 = ~n470 & ~n667;
  assign n790 = ~n403 & ~n513;
  assign n791 = n98 & n106;
  assign n792 = ~n168 & ~n791;
  assign n793 = ~n161 & ~n245;
  assign n794 = n792 & n793;
  assign n795 = n790 & n794;
  assign n796 = n789 & n795;
  assign n797 = n622 & n796;
  assign n798 = ~n177 & n797;
  assign n799 = ~n396 & n798;
  assign n800 = ~n277 & n799;
  assign n801 = n788 & n800;
  assign n802 = ~n449 & n801;
  assign n803 = n96 & n114;
  assign n804 = ~n326 & ~n511;
  assign n805 = ~n495 & ~n514;
  assign n806 = ~n296 & ~n492;
  assign n807 = ~n422 & n806;
  assign n808 = ~n375 & n807;
  assign n809 = n113 & n174;
  assign n810 = ~n430 & ~n809;
  assign n811 = ~n150 & ~n284;
  assign n812 = ~n149 & ~n417;
  assign n813 = ~n623 & ~n641;
  assign n814 = ~n666 & n813;
  assign n815 = ~n169 & ~n620;
  assign n816 = ~n672 & n815;
  assign n817 = n814 & n816;
  assign n818 = n812 & n817;
  assign n819 = n811 & n818;
  assign n820 = n810 & n819;
  assign n821 = ~n228 & n820;
  assign n822 = ~n243 & n821;
  assign n823 = ~n366 & n822;
  assign n824 = ~n562 & n823;
  assign n825 = n90 & n176;
  assign n826 = ~n246 & ~n420;
  assign n827 = ~n295 & ~n564;
  assign n828 = n826 & n827;
  assign n829 = ~n121 & n828;
  assign n830 = ~n825 & n829;
  assign n831 = ~n504 & ~n518;
  assign n832 = ~n270 & n831;
  assign n833 = n467 & n832;
  assign n834 = n830 & n833;
  assign n835 = n824 & n834;
  assign n836 = n808 & n835;
  assign n837 = n805 & n836;
  assign n838 = n804 & n837;
  assign n839 = ~n509 & n838;
  assign n840 = ~n557 & n839;
  assign n841 = ~n254 & n840;
  assign n842 = ~n803 & n841;
  assign n843 = ~n280 & n842;
  assign n844 = ~n532 & n843;
  assign n845 = n120 & n654;
  assign n846 = ~n189 & n845;
  assign n847 = n88 & n153;
  assign n848 = ~n558 & ~n847;
  assign n849 = ~n223 & n848;
  assign n850 = ~n617 & n849;
  assign n851 = ~n353 & n850;
  assign n852 = n846 & n851;
  assign n853 = n844 & n852;
  assign n854 = n802 & n853;
  assign n855 = n787 & n854;
  assign n856 = n772 & n855;
  assign n857 = n770 & n856;
  assign n858 = ~n713 & n857;
  assign n859 = ~n151 & n858;
  assign n860 = ~n299 & n859;
  assign n861 = ~n639 & n860;
  assign n862 = ~n496 & n861;
  assign n863 = ~n142 & n862;
  assign n864 = ~n468 & n863;
  assign n865 = ~n712 & n864;
  assign n866 = ~n489 & n865;
  assign n867 = ~n188 & n866;
  assign n868 = ~n710 & ~n867;
  assign n869 = ~n224 & ~n243;
  assign n870 = ~n155 & ~n254;
  assign n871 = ~n777 & n870;
  assign n872 = ~n304 & n871;
  assign n873 = ~n144 & ~n713;
  assign n874 = ~n236 & ~n272;
  assign n875 = n80 & n96;
  assign n876 = ~n301 & ~n513;
  assign n877 = ~n330 & ~n715;
  assign n878 = n876 & n877;
  assign n879 = ~n602 & n878;
  assign n880 = ~n205 & n879;
  assign n881 = ~n325 & n880;
  assign n882 = ~n875 & n881;
  assign n883 = n78 & n83;
  assign n884 = n106 & n117;
  assign n885 = ~n86 & ~n296;
  assign n886 = n83 & n113;
  assign n887 = ~n426 & ~n562;
  assign n888 = ~n326 & ~n637;
  assign n889 = ~n496 & n888;
  assign n890 = n887 & n889;
  assign n891 = ~n594 & n890;
  assign n892 = ~n419 & n891;
  assign n893 = ~n417 & n892;
  assign n894 = ~n886 & n893;
  assign n895 = ~n429 & n894;
  assign n896 = ~n425 & ~n489;
  assign n897 = ~n338 & ~n427;
  assign n898 = ~n354 & n719;
  assign n899 = ~n393 & n898;
  assign n900 = n897 & n899;
  assign n901 = n851 & n900;
  assign n902 = n539 & n901;
  assign n903 = n128 & n902;
  assign n904 = n896 & n903;
  assign n905 = n399 & n904;
  assign n906 = n895 & n905;
  assign n907 = n507 & n906;
  assign n908 = n885 & n907;
  assign n909 = ~n229 & n908;
  assign n910 = n572 & n909;
  assign n911 = ~n619 & n910;
  assign n912 = ~n884 & n911;
  assign n913 = ~n825 & n912;
  assign n914 = ~n331 & n913;
  assign n915 = ~n883 & n914;
  assign n916 = ~n428 & n915;
  assign n917 = ~n242 & ~n335;
  assign n918 = ~n771 & n917;
  assign n919 = ~n194 & ~n589;
  assign n920 = ~n130 & n919;
  assign n921 = ~n633 & n920;
  assign n922 = n179 & n921;
  assign n923 = n918 & n922;
  assign n924 = ~n255 & n923;
  assign n925 = ~n189 & n924;
  assign n926 = ~n328 & n925;
  assign n927 = ~n809 & n926;
  assign n928 = ~n461 & n927;
  assign n929 = ~n395 & n928;
  assign n930 = ~n145 & n929;
  assign n931 = ~n251 & n930;
  assign n932 = n88 & n129;
  assign n933 = ~n436 & ~n932;
  assign n934 = n235 & n933;
  assign n935 = n454 & n934;
  assign n936 = ~n142 & n935;
  assign n937 = ~n119 & ~n438;
  assign n938 = ~n281 & n937;
  assign n939 = ~n352 & n938;
  assign n940 = ~n623 & n939;
  assign n941 = ~n147 & ~n295;
  assign n942 = n475 & n941;
  assign n943 = n940 & n942;
  assign n944 = n936 & n943;
  assign n945 = n931 & n944;
  assign n946 = n916 & n945;
  assign n947 = n882 & n946;
  assign n948 = n874 & n947;
  assign n949 = n873 & n948;
  assign n950 = n872 & n949;
  assign n951 = n423 & n950;
  assign n952 = n869 & n951;
  assign n953 = ~n746 & n952;
  assign n954 = ~n355 & n953;
  assign n955 = ~n400 & n954;
  assign n956 = ~n374 & n955;
  assign n957 = ~n492 & n956;
  assign n958 = ~n158 & n957;
  assign n959 = ~n867 & ~n958;
  assign n960 = ~n111 & ~n254;
  assign n961 = n94 & n98;
  assign n962 = ~n397 & ~n961;
  assign n963 = n960 & n962;
  assign n964 = ~n352 & n963;
  assign n965 = ~n884 & n964;
  assign n966 = ~n102 & n965;
  assign n967 = ~n240 & n966;
  assign n968 = ~n81 & ~n337;
  assign n969 = ~n276 & n968;
  assign n970 = ~n299 & n969;
  assign n971 = ~n513 & n970;
  assign n972 = ~n165 & n971;
  assign n973 = ~n791 & n972;
  assign n974 = ~n531 & n973;
  assign n975 = ~n489 & n974;
  assign n976 = ~n883 & n975;
  assign n977 = ~n394 & ~n429;
  assign n978 = ~n326 & ~n639;
  assign n979 = ~n353 & ~n620;
  assign n980 = n106 & n166;
  assign n981 = ~n203 & ~n286;
  assign n982 = ~n366 & n981;
  assign n983 = n515 & n982;
  assign n984 = ~n339 & n983;
  assign n985 = ~n118 & n984;
  assign n986 = ~n980 & n985;
  assign n987 = ~n192 & n986;
  assign n988 = ~n173 & n987;
  assign n989 = ~n436 & ~n589;
  assign n990 = ~n466 & ~n493;
  assign n991 = ~n149 & ~n617;
  assign n992 = ~n825 & n991;
  assign n993 = n990 & n992;
  assign n994 = n989 & n993;
  assign n995 = n988 & n994;
  assign n996 = n510 & n995;
  assign n997 = n294 & n996;
  assign n998 = n238 & n997;
  assign n999 = n979 & n998;
  assign n1000 = n978 & n999;
  assign n1001 = n227 & n1000;
  assign n1002 = n418 & n1001;
  assign n1003 = ~n746 & n1002;
  assign n1004 = ~n177 & n1003;
  assign n1005 = ~n689 & n1004;
  assign n1006 = ~n164 & n1005;
  assign n1007 = ~n338 & n1006;
  assign n1008 = ~n125 & n1007;
  assign n1009 = ~n150 & ~n252;
  assign n1010 = n131 & n160;
  assign n1011 = n113 & n153;
  assign n1012 = ~n400 & ~n672;
  assign n1013 = ~n427 & n1012;
  assign n1014 = ~n1011 & n1013;
  assign n1015 = ~n435 & n1014;
  assign n1016 = ~n932 & n1015;
  assign n1017 = ~n130 & n1016;
  assign n1018 = ~n623 & n1017;
  assign n1019 = ~n1010 & n1018;
  assign n1020 = ~n564 & n1019;
  assign n1021 = ~n190 & ~n224;
  assign n1022 = ~n233 & n1021;
  assign n1023 = ~n490 & n1022;
  assign n1024 = ~n249 & n1023;
  assign n1025 = ~n154 & ~n273;
  assign n1026 = n405 & n1025;
  assign n1027 = n1024 & n1026;
  assign n1028 = n1020 & n1027;
  assign n1029 = n431 & ~n803;
  assign n1030 = n1028 & n1029;
  assign n1031 = n244 & n1030;
  assign n1032 = n1009 & n1031;
  assign n1033 = n747 & n1032;
  assign n1034 = ~n123 & n1033;
  assign n1035 = ~n426 & n1034;
  assign n1036 = ~n416 & n1035;
  assign n1037 = ~n142 & n1036;
  assign n1038 = ~n422 & n1037;
  assign n1039 = ~n251 & n1038;
  assign n1040 = ~n304 & ~n557;
  assign n1041 = n570 & n1040;
  assign n1042 = ~n847 & n1041;
  assign n1043 = ~n152 & n1042;
  assign n1044 = ~n171 & n1043;
  assign n1045 = ~n136 & n282;
  assign n1046 = ~n167 & ~n246;
  assign n1047 = ~n163 & n1046;
  assign n1048 = n1045 & n1047;
  assign n1049 = n1044 & n1048;
  assign n1050 = n1039 & n1049;
  assign n1051 = n1008 & n1050;
  assign n1052 = n977 & n1051;
  assign n1053 = n622 & n1052;
  assign n1054 = n976 & n1053;
  assign n1055 = n967 & n1054;
  assign n1056 = n885 & n1055;
  assign n1057 = ~n602 & n1056;
  assign n1058 = ~n506 & n1057;
  assign n1059 = ~n425 & n1058;
  assign n1060 = ~n157 & n1059;
  assign n1061 = ~n958 & ~n1060;
  assign n1062 = n131 & n174;
  assign n1063 = ~n177 & ~n416;
  assign n1064 = ~n419 & ~n1011;
  assign n1065 = ~n337 & n1064;
  assign n1066 = ~n398 & n1065;
  assign n1067 = ~n400 & n1066;
  assign n1068 = ~n167 & n1067;
  assign n1069 = ~n875 & n1068;
  assign n1070 = ~n252 & ~n509;
  assign n1071 = ~n165 & ~n237;
  assign n1072 = n110 & n124;
  assign n1073 = ~n155 & ~n1072;
  assign n1074 = n1071 & n1073;
  assign n1075 = n1070 & n1074;
  assign n1076 = ~n301 & n1075;
  assign n1077 = ~n641 & n1076;
  assign n1078 = ~n149 & n1077;
  assign n1079 = ~n107 & n1078;
  assign n1080 = ~n173 & n1079;
  assign n1081 = ~n189 & ~n296;
  assign n1082 = ~n537 & n1081;
  assign n1083 = ~n422 & n1082;
  assign n1084 = ~n451 & n1083;
  assign n1085 = ~n274 & ~n531;
  assign n1086 = n256 & n1085;
  assign n1087 = n1084 & n1086;
  assign n1088 = n1080 & n1087;
  assign n1089 = n1069 & n1088;
  assign n1090 = n1063 & n1089;
  assign n1091 = n159 & n1090;
  assign n1092 = n570 & n1091;
  assign n1093 = ~n115 & n1092;
  assign n1094 = ~n1062 & n1093;
  assign n1095 = ~n298 & n1094;
  assign n1096 = ~n589 & n1095;
  assign n1097 = ~n366 & n1096;
  assign n1098 = ~n340 & n1097;
  assign n1099 = ~n371 & n1098;
  assign n1100 = ~n271 & n1099;
  assign n1101 = n148 & n174;
  assign n1102 = n85 & n114;
  assign n1103 = ~n466 & ~n1102;
  assign n1104 = n122 & n199;
  assign n1105 = ~n519 & ~n1104;
  assign n1106 = ~n603 & n1105;
  assign n1107 = ~n771 & n1106;
  assign n1108 = ~n171 & ~n752;
  assign n1109 = ~n712 & n1108;
  assign n1110 = n1107 & n1109;
  assign n1111 = n1103 & n1110;
  assign n1112 = ~n136 & n1111;
  assign n1113 = ~n397 & n1112;
  assign n1114 = ~n462 & n1113;
  assign n1115 = ~n847 & n1114;
  assign n1116 = ~n1101 & n1115;
  assign n1117 = ~n435 & n1116;
  assign n1118 = ~n395 & n1117;
  assign n1119 = ~n127 & n1118;
  assign n1120 = ~n239 & ~n246;
  assign n1121 = ~n273 & n1120;
  assign n1122 = ~n402 & n1121;
  assign n1123 = ~n716 & n1122;
  assign n1124 = ~n144 & n1123;
  assign n1125 = ~n201 & n1124;
  assign n1126 = ~n332 & n1125;
  assign n1127 = n126 & n160;
  assign n1128 = ~n883 & ~n1127;
  assign n1129 = ~n428 & ~n469;
  assign n1130 = ~n151 & ~n557;
  assign n1131 = ~n506 & n1130;
  assign n1132 = ~n424 & ~n803;
  assign n1133 = ~n121 & ~n276;
  assign n1134 = ~n490 & n1133;
  assign n1135 = ~n666 & n1134;
  assign n1136 = ~n299 & ~n426;
  assign n1137 = ~n673 & n1136;
  assign n1138 = ~n394 & n1137;
  assign n1139 = ~n205 & ~n292;
  assign n1140 = ~n564 & n1139;
  assign n1141 = ~n270 & ~n338;
  assign n1142 = ~n275 & n1141;
  assign n1143 = ~n163 & n1142;
  assign n1144 = n1140 & n1143;
  assign n1145 = n1138 & n1144;
  assign n1146 = n1135 & n1145;
  assign n1147 = n1132 & n1146;
  assign n1148 = n936 & n1147;
  assign n1149 = n1131 & n1148;
  assign n1150 = n1129 & n1149;
  assign n1151 = n654 & n1150;
  assign n1152 = n1128 & n1151;
  assign n1153 = ~n637 & n1152;
  assign n1154 = ~n367 & n1153;
  assign n1155 = ~n304 & ~n1010;
  assign n1156 = n773 & n979;
  assign n1157 = ~n132 & n1156;
  assign n1158 = ~n655 & n1157;
  assign n1159 = ~n99 & ~n305;
  assign n1160 = ~n293 & n1159;
  assign n1161 = ~n191 & ~n468;
  assign n1162 = ~n281 & n1161;
  assign n1163 = ~n714 & n1162;
  assign n1164 = n1160 & n1163;
  assign n1165 = n776 & n1164;
  assign n1166 = n1158 & n1165;
  assign n1167 = n1155 & n1166;
  assign n1168 = n1154 & n1167;
  assign n1169 = n1126 & n1168;
  assign n1170 = n1119 & n1169;
  assign n1171 = n665 & n1170;
  assign n1172 = n1100 & n1171;
  assign n1173 = n896 & n1172;
  assign n1174 = n937 & n1173;
  assign n1175 = ~n617 & n1174;
  assign n1176 = ~n495 & n1175;
  assign n1177 = ~n460 & n1176;
  assign n1178 = ~n562 & n1177;
  assign n1179 = ~n1060 & ~n1178;
  assign n1180 = ~n135 & ~n657;
  assign n1181 = ~n152 & ~n505;
  assign n1182 = ~n81 & ~n329;
  assign n1183 = ~n419 & ~n435;
  assign n1184 = n238 & n937;
  assign n1185 = ~n194 & n1184;
  assign n1186 = n675 & n1185;
  assign n1187 = n751 & n1186;
  assign n1188 = n1155 & n1187;
  assign n1189 = n787 & n1188;
  assign n1190 = n1183 & n1189;
  assign n1191 = n1182 & n1190;
  assign n1192 = ~n301 & n1191;
  assign n1193 = ~n136 & n1192;
  assign n1194 = ~n111 & n1193;
  assign n1195 = ~n354 & n1194;
  assign n1196 = ~n224 & n1195;
  assign n1197 = ~n884 & n1196;
  assign n1198 = ~n173 & n1197;
  assign n1199 = ~n164 & n1198;
  assign n1200 = ~n536 & n1199;
  assign n1201 = ~n603 & n1200;
  assign n1202 = ~n655 & n1201;
  assign n1203 = n122 & n129;
  assign n1204 = ~n569 & ~n980;
  assign n1205 = ~n340 & ~n527;
  assign n1206 = ~n875 & n1205;
  assign n1207 = n1204 & n1206;
  assign n1208 = ~n327 & n1207;
  assign n1209 = ~n228 & n1208;
  assign n1210 = ~n1203 & n1209;
  assign n1211 = ~n325 & n1210;
  assign n1212 = ~n154 & ~n254;
  assign n1213 = ~n400 & n1212;
  assign n1214 = ~n102 & n1213;
  assign n1215 = ~n331 & n1214;
  assign n1216 = ~n589 & n1215;
  assign n1217 = ~n167 & ~n563;
  assign n1218 = ~n306 & n1217;
  assign n1219 = ~n251 & n1218;
  assign n1220 = ~n422 & ~n656;
  assign n1221 = ~n222 & n1220;
  assign n1222 = n982 & n1221;
  assign n1223 = n1219 & n1222;
  assign n1224 = n1216 & n1223;
  assign n1225 = n1154 & n1224;
  assign n1226 = n802 & n1225;
  assign n1227 = n1211 & n1226;
  assign n1228 = n1202 & n1227;
  assign n1229 = n1181 & n1228;
  assign n1230 = n1180 & n1229;
  assign n1231 = ~n518 & n1230;
  assign n1232 = ~n374 & n1231;
  assign n1233 = ~n601 & n1232;
  assign n1234 = ~n200 & n1233;
  assign n1235 = ~n295 & n1234;
  assign n1236 = ~n1178 & ~n1235;
  assign n1237 = ~n224 & ~n397;
  assign n1238 = ~n150 & ~n417;
  assign n1239 = ~n305 & n1238;
  assign n1240 = ~n374 & n1239;
  assign n1241 = n590 & n1240;
  assign n1242 = ~n402 & n1241;
  assign n1243 = ~n496 & n1242;
  assign n1244 = ~n424 & n1243;
  assign n1245 = ~n277 & n1244;
  assign n1246 = n153 & n269;
  assign n1247 = ~n274 & ~n469;
  assign n1248 = ~n352 & ~n1101;
  assign n1249 = ~n192 & ~n251;
  assign n1250 = n303 & n1249;
  assign n1251 = ~n673 & n1250;
  assign n1252 = ~n371 & ~n504;
  assign n1253 = ~n368 & ~n771;
  assign n1254 = ~n255 & ~n562;
  assign n1255 = ~n99 & ~n249;
  assign n1256 = n814 & n1255;
  assign n1257 = n734 & n1256;
  assign n1258 = n1254 & n1257;
  assign n1259 = n1253 & n1258;
  assign n1260 = n1252 & n1259;
  assign n1261 = ~n495 & n1260;
  assign n1262 = ~n296 & n1261;
  assign n1263 = ~n961 & n1262;
  assign n1264 = ~n567 & n1263;
  assign n1265 = n244 & ~n980;
  assign n1266 = ~n537 & n1265;
  assign n1267 = ~n170 & n1266;
  assign n1268 = ~n86 & n1267;
  assign n1269 = ~n427 & ~n449;
  assign n1270 = ~n329 & n1269;
  assign n1271 = ~n884 & n1270;
  assign n1272 = ~n154 & ~n514;
  assign n1273 = n533 & ~n617;
  assign n1274 = ~n398 & n1273;
  assign n1275 = n1272 & n1274;
  assign n1276 = n1271 & n1275;
  assign n1277 = n1103 & n1276;
  assign n1278 = n1268 & n1277;
  assign n1279 = n1264 & n1278;
  assign n1280 = n1251 & n1279;
  assign n1281 = n235 & n1280;
  assign n1282 = n285 & n1281;
  assign n1283 = n1248 & n1282;
  assign n1284 = n1247 & n1283;
  assign n1285 = ~n1246 & n1284;
  assign n1286 = ~n426 & n1285;
  assign n1287 = ~n189 & n1286;
  assign n1288 = ~n460 & n1287;
  assign n1289 = ~n287 & n1288;
  assign n1290 = ~n932 & n1289;
  assign n1291 = ~n569 & n1290;
  assign n1292 = ~n558 & ~n803;
  assign n1293 = ~n375 & ~n639;
  assign n1294 = ~n273 & n1293;
  assign n1295 = n735 & n1294;
  assign n1296 = n359 & n1295;
  assign n1297 = ~n509 & n1296;
  assign n1298 = ~n190 & n1297;
  assign n1299 = ~n461 & n1298;
  assign n1300 = ~n601 & n1299;
  assign n1301 = ~n191 & n1300;
  assign n1302 = ~n436 & n1301;
  assign n1303 = ~n125 & n1302;
  assign n1304 = ~n81 & n1303;
  assign n1305 = ~n633 & n1304;
  assign n1306 = n78 & n110;
  assign n1307 = ~n395 & ~n689;
  assign n1308 = ~n453 & n1307;
  assign n1309 = ~n1306 & n1308;
  assign n1310 = ~n619 & n1309;
  assign n1311 = ~n290 & n1310;
  assign n1312 = ~n331 & n1311;
  assign n1313 = ~n270 & n1312;
  assign n1314 = ~n394 & ~n396;
  assign n1315 = ~n451 & n1314;
  assign n1316 = n1139 & n1315;
  assign n1317 = ~n330 & n1316;
  assign n1318 = ~n339 & n1317;
  assign n1319 = ~n146 & n1318;
  assign n1320 = ~n492 & n1319;
  assign n1321 = ~n714 & n1320;
  assign n1322 = ~n304 & n1321;
  assign n1323 = ~n337 & n1322;
  assign n1324 = ~n518 & ~n568;
  assign n1325 = ~n157 & n1324;
  assign n1326 = ~n470 & n1325;
  assign n1327 = ~n657 & n1326;
  assign n1328 = ~n428 & n1327;
  assign n1329 = ~n149 & ~n602;
  assign n1330 = ~n847 & ~n886;
  assign n1331 = ~n237 & n1330;
  assign n1332 = ~n200 & ~n299;
  assign n1333 = ~n161 & n1332;
  assign n1334 = n1331 & n1333;
  assign n1335 = n1329 & n1334;
  assign n1336 = n1328 & n1335;
  assign n1337 = n1323 & n1336;
  assign n1338 = n731 & n1337;
  assign n1339 = n1313 & n1338;
  assign n1340 = ~n746 & n1339;
  assign n1341 = ~n281 & n1340;
  assign n1342 = ~n335 & n1341;
  assign n1343 = ~n115 & n1342;
  assign n1344 = ~n239 & n1343;
  assign n1345 = ~n226 & n1344;
  assign n1346 = ~n118 & ~n354;
  assign n1347 = ~n367 & ~n400;
  assign n1348 = n1346 & n1347;
  assign n1349 = n830 & n1348;
  assign n1350 = n1345 & n1349;
  assign n1351 = n1305 & n1350;
  assign n1352 = n1292 & n1351;
  assign n1353 = n1291 & n1352;
  assign n1354 = n1245 & n1353;
  assign n1355 = n937 & n1354;
  assign n1356 = n1237 & n1355;
  assign n1357 = ~n194 & n1356;
  assign n1358 = ~n328 & n1357;
  assign n1359 = ~n175 & n1358;
  assign n1360 = ~n637 & n1359;
  assign n1361 = ~n422 & n1360;
  assign n1362 = ~n468 & n1361;
  assign n1363 = ~n531 & n1362;
  assign n1364 = ~n366 & n1363;
  assign n1365 = ~n1235 & ~n1364;
  assign n1366 = ~n225 & ~n601;
  assign n1367 = ~n170 & ~n273;
  assign n1368 = ~n191 & ~n352;
  assign n1369 = ~n272 & n1368;
  assign n1370 = ~n305 & ~n506;
  assign n1371 = ~n246 & n1370;
  assign n1372 = ~n712 & n1371;
  assign n1373 = n1369 & n1372;
  assign n1374 = n1367 & n1373;
  assign n1375 = ~n111 & n1374;
  assign n1376 = ~n147 & n1375;
  assign n1377 = ~n884 & n1376;
  assign n1378 = ~n302 & n1377;
  assign n1379 = ~n531 & ~n1306;
  assign n1380 = ~n329 & ~n474;
  assign n1381 = ~n229 & n1380;
  assign n1382 = ~n354 & n1381;
  assign n1383 = ~n296 & n1382;
  assign n1384 = ~n589 & n1383;
  assign n1385 = ~n330 & ~n803;
  assign n1386 = ~n791 & n1385;
  assign n1387 = ~n372 & n1386;
  assign n1388 = ~n331 & ~n932;
  assign n1389 = ~n203 & ~n461;
  assign n1390 = ~n620 & n1389;
  assign n1391 = ~n519 & n1390;
  assign n1392 = ~n275 & ~n375;
  assign n1393 = ~n403 & ~n1102;
  assign n1394 = ~n200 & n1393;
  assign n1395 = n1392 & n1394;
  assign n1396 = n846 & n1395;
  assign n1397 = n1391 & n1396;
  assign n1398 = n1388 & n1397;
  assign n1399 = n1387 & n1398;
  assign n1400 = n1384 & n1399;
  assign n1401 = n1379 & n1400;
  assign n1402 = n1180 & n1401;
  assign n1403 = n1128 & n1402;
  assign n1404 = ~n462 & n1403;
  assign n1405 = ~n232 & n1404;
  assign n1406 = ~n223 & n1405;
  assign n1407 = ~n623 & n1406;
  assign n1408 = ~n107 & ~n715;
  assign n1409 = ~n633 & ~n961;
  assign n1410 = n1408 & n1409;
  assign n1411 = n789 & n1410;
  assign n1412 = ~n752 & n1411;
  assign n1413 = ~n278 & n1412;
  assign n1414 = ~n326 & n1413;
  assign n1415 = ~n490 & n1414;
  assign n1416 = ~n145 & n1415;
  assign n1417 = ~n99 & n1416;
  assign n1418 = ~n672 & n1417;
  assign n1419 = ~n271 & n1418;
  assign n1420 = ~n367 & ~n496;
  assign n1421 = ~n673 & n1420;
  assign n1422 = ~n86 & n1421;
  assign n1423 = ~n91 & ~n164;
  assign n1424 = ~n165 & ~n495;
  assign n1425 = ~n619 & ~n771;
  assign n1426 = ~n276 & ~n592;
  assign n1427 = ~n689 & n1426;
  assign n1428 = ~n429 & n1427;
  assign n1429 = n1425 & n1428;
  assign n1430 = n1219 & n1429;
  assign n1431 = n1424 & n1430;
  assign n1432 = n1063 & n1431;
  assign n1433 = ~n527 & n1432;
  assign n1434 = ~n102 & n1433;
  assign n1435 = ~n231 & n1434;
  assign n1436 = ~n395 & ~n571;
  assign n1437 = ~n825 & n1436;
  assign n1438 = ~n289 & ~n1062;
  assign n1439 = ~n602 & ~n641;
  assign n1440 = ~n150 & n1439;
  assign n1441 = n1065 & n1440;
  assign n1442 = n1438 & n1441;
  assign n1443 = n1437 & n1442;
  assign n1444 = n604 & n1443;
  assign n1445 = n1435 & n1444;
  assign n1446 = n1139 & n1445;
  assign n1447 = n896 & n1446;
  assign n1448 = n827 & n1447;
  assign n1449 = n1237 & n1448;
  assign n1450 = ~n847 & n1449;
  assign n1451 = ~n417 & n1450;
  assign n1452 = ~n228 & n1451;
  assign n1453 = ~n173 & n1452;
  assign n1454 = ~n95 & n1453;
  assign n1455 = n454 & n1454;
  assign n1456 = ~n639 & n1455;
  assign n1457 = ~n152 & ~n567;
  assign n1458 = ~n161 & n1457;
  assign n1459 = n1456 & n1458;
  assign n1460 = n1423 & n1459;
  assign n1461 = n1422 & n1460;
  assign n1462 = n1419 & n1461;
  assign n1463 = n1407 & n1462;
  assign n1464 = n1378 & n1463;
  assign n1465 = n1366 & n1464;
  assign n1466 = n1269 & n1465;
  assign n1467 = ~n558 & n1466;
  assign n1468 = ~n509 & n1467;
  assign n1469 = ~n149 & n1468;
  assign n1470 = ~n402 & n1469;
  assign n1471 = ~n777 & n1470;
  assign n1472 = ~n132 & n1471;
  assign n1473 = ~n1364 & ~n1472;
  assign n1474 = ~n427 & ~n568;
  assign n1475 = ~n283 & n1474;
  assign n1476 = ~n232 & ~n332;
  assign n1477 = ~n395 & ~n416;
  assign n1478 = ~n374 & n1477;
  assign n1479 = ~n496 & ~n746;
  assign n1480 = ~n249 & ~n655;
  assign n1481 = n253 & n1384;
  assign n1482 = ~n284 & n1481;
  assign n1483 = ~n715 & n1482;
  assign n1484 = ~n394 & n1483;
  assign n1485 = ~n132 & n1484;
  assign n1486 = ~n470 & n1485;
  assign n1487 = ~n1010 & n1486;
  assign n1488 = ~n158 & n1487;
  assign n1489 = ~n107 & ~n1011;
  assign n1490 = ~n170 & n1489;
  assign n1491 = ~n435 & n1490;
  assign n1492 = ~n884 & n1491;
  assign n1493 = ~n331 & n1492;
  assign n1494 = ~n157 & n1493;
  assign n1495 = ~n295 & n1494;
  assign n1496 = ~n127 & n1495;
  assign n1497 = ~n155 & ~n809;
  assign n1498 = ~n513 & ~n752;
  assign n1499 = ~n425 & n1498;
  assign n1500 = n1497 & n1499;
  assign n1501 = n1496 & n1500;
  assign n1502 = n1488 & n1501;
  assign n1503 = n1480 & n1502;
  assign n1504 = n1479 & n1503;
  assign n1505 = n1478 & n1504;
  assign n1506 = ~n602 & n1505;
  assign n1507 = ~n334 & n1506;
  assign n1508 = ~n173 & n1507;
  assign n1509 = ~n657 & n1508;
  assign n1510 = ~n569 & n1509;
  assign n1511 = ~n270 & n1510;
  assign n1512 = ~n364 & n960;
  assign n1513 = ~n123 & n1512;
  assign n1514 = ~n713 & n1513;
  assign n1515 = ~n327 & n1514;
  assign n1516 = ~n177 & n1515;
  assign n1517 = ~n275 & n1516;
  assign n1518 = ~n825 & n1517;
  assign n1519 = ~n240 & n1518;
  assign n1520 = ~n272 & n1519;
  assign n1521 = ~n771 & n1520;
  assign n1522 = ~n223 & ~n562;
  assign n1523 = ~n149 & ~n298;
  assign n1524 = ~n146 & ~n495;
  assign n1525 = ~n167 & n1524;
  assign n1526 = ~n603 & n1525;
  assign n1527 = ~n489 & n1526;
  assign n1528 = ~n353 & ~n396;
  assign n1529 = ~n326 & n1528;
  assign n1530 = ~n449 & n1529;
  assign n1531 = ~n293 & ~n666;
  assign n1532 = n1129 & n1531;
  assign n1533 = ~n716 & n1532;
  assign n1534 = n1331 & n1533;
  assign n1535 = n1530 & n1534;
  assign n1536 = n723 & n1535;
  assign n1537 = n439 & n1536;
  assign n1538 = n1527 & n1537;
  assign n1539 = n1105 & n1538;
  assign n1540 = n1305 & n1539;
  assign n1541 = n1523 & n1540;
  assign n1542 = n1426 & n1541;
  assign n1543 = n590 & n1542;
  assign n1544 = n1522 & n1543;
  assign n1545 = ~n339 & n1544;
  assign n1546 = ~n505 & n1545;
  assign n1547 = ~n306 & n1546;
  assign n1548 = ~n304 & n1547;
  assign n1549 = ~n525 & n1548;
  assign n1550 = ~n274 & ~n558;
  assign n1551 = n202 & n282;
  assign n1552 = n1550 & n1551;
  assign n1553 = ~n980 & n1552;
  assign n1554 = ~n453 & n1553;
  assign n1555 = ~n277 & n1554;
  assign n1556 = ~n130 & ~n366;
  assign n1557 = ~n271 & ~n462;
  assign n1558 = n1556 & n1557;
  assign n1559 = n1555 & n1558;
  assign n1560 = n1549 & n1559;
  assign n1561 = n1521 & n1560;
  assign n1562 = n631 & n1561;
  assign n1563 = n1511 & n1562;
  assign n1564 = n1476 & n1563;
  assign n1565 = n1475 & n1564;
  assign n1566 = n288 & n1565;
  assign n1567 = n1379 & n1566;
  assign n1568 = ~n424 & n1567;
  assign n1569 = ~n205 & n1568;
  assign n1570 = ~n537 & n1569;
  assign n1571 = ~n161 & n1570;
  assign n1572 = ~n429 & n1571;
  assign n1573 = ~n1472 & ~n1572;
  assign n1574 = ~n284 & ~n532;
  assign n1575 = ~n170 & ~n328;
  assign n1576 = ~n142 & ~n714;
  assign n1577 = ~n272 & ~n1203;
  assign n1578 = ~n452 & n772;
  assign n1579 = n1577 & n1578;
  assign n1580 = n1181 & n1579;
  assign n1581 = n873 & n1580;
  assign n1582 = n235 & n1581;
  assign n1583 = ~n617 & n1582;
  assign n1584 = ~n275 & n1583;
  assign n1585 = ~n86 & n1584;
  assign n1586 = ~n639 & ~n657;
  assign n1587 = ~n274 & ~n504;
  assign n1588 = ~n201 & n1587;
  assign n1589 = n1428 & n1588;
  assign n1590 = n1586 & n1589;
  assign n1591 = n1585 & n1590;
  assign n1592 = n1480 & n1591;
  assign n1593 = n120 & n1592;
  assign n1594 = n1576 & n1593;
  assign n1595 = n731 & n1594;
  assign n1596 = n156 & n1595;
  assign n1597 = ~n254 & n1596;
  assign n1598 = ~n641 & n1597;
  assign n1599 = ~n171 & n1598;
  assign n1600 = ~n287 & n1599;
  assign n1601 = ~n177 & ~n236;
  assign n1602 = ~n161 & ~n354;
  assign n1603 = ~n190 & ~n280;
  assign n1604 = ~n603 & ~n1011;
  assign n1605 = n1603 & n1604;
  assign n1606 = n294 & n1605;
  assign n1607 = ~n400 & n1606;
  assign n1608 = ~n102 & n1607;
  assign n1609 = ~n496 & n1608;
  assign n1610 = ~n246 & n1609;
  assign n1611 = ~n492 & ~n1010;
  assign n1612 = ~n1246 & n1611;
  assign n1613 = ~n327 & n1612;
  assign n1614 = ~n637 & n1613;
  assign n1615 = ~n438 & n1614;
  assign n1616 = ~n111 & ~n601;
  assign n1617 = ~n672 & n1616;
  assign n1618 = ~n329 & ~n620;
  assign n1619 = ~n980 & n1618;
  assign n1620 = ~n337 & n1619;
  assign n1621 = ~n449 & n1620;
  assign n1622 = n1617 & n1621;
  assign n1623 = n1615 & n1622;
  assign n1624 = n1610 & n1623;
  assign n1625 = n1602 & n1624;
  assign n1626 = ~n301 & n1625;
  assign n1627 = ~n558 & n1626;
  assign n1628 = ~n461 & n1627;
  assign n1629 = ~n91 & n1628;
  assign n1630 = ~n416 & n1629;
  assign n1631 = ~n368 & n1630;
  assign n1632 = ~n468 & n1631;
  assign n1633 = ~n623 & n1632;
  assign n1634 = ~n277 & n1633;
  assign n1635 = ~n489 & n1634;
  assign n1636 = ~n424 & ~n1306;
  assign n1637 = ~n278 & n1636;
  assign n1638 = ~n619 & n1637;
  assign n1639 = ~n374 & n1638;
  assign n1640 = ~n251 & n1639;
  assign n1641 = ~n339 & ~n427;
  assign n1642 = ~n273 & n1641;
  assign n1643 = ~n712 & n1642;
  assign n1644 = ~n228 & ~n777;
  assign n1645 = ~n223 & n1254;
  assign n1646 = ~n331 & n1645;
  assign n1647 = n1644 & n1646;
  assign n1648 = n1643 & n1647;
  assign n1649 = n1640 & n1648;
  assign n1650 = n1635 & n1649;
  assign n1651 = n1601 & n1650;
  assign n1652 = n1600 & n1651;
  assign n1653 = n1575 & n1652;
  assign n1654 = n423 & n1653;
  assign n1655 = n745 & n1654;
  assign n1656 = n1248 & n1655;
  assign n1657 = n1574 & n1656;
  assign n1658 = n359 & n1657;
  assign n1659 = ~n151 & n1658;
  assign n1660 = ~n326 & n1659;
  assign n1661 = ~n568 & n1660;
  assign n1662 = ~n286 & n1661;
  assign n1663 = ~n567 & n1662;
  assign n1664 = ~n1104 & n1663;
  assign n1665 = ~n271 & n1664;
  assign n1666 = ~n1572 & ~n1665;
  assign n1667 = ~n132 & ~n249;
  assign n1668 = ~n91 & ~n462;
  assign n1669 = ~n428 & n788;
  assign n1670 = n849 & n1669;
  assign n1671 = n933 & n1670;
  assign n1672 = n1475 & n1671;
  assign n1673 = n1668 & n1672;
  assign n1674 = ~n111 & n1673;
  assign n1675 = ~n716 & n1674;
  assign n1676 = ~n425 & n1675;
  assign n1677 = ~n589 & n1676;
  assign n1678 = ~n531 & n1677;
  assign n1679 = ~n231 & n1678;
  assign n1680 = ~n714 & ~n1104;
  assign n1681 = ~n633 & n1680;
  assign n1682 = n303 & n1681;
  assign n1683 = n790 & n1682;
  assign n1684 = ~n364 & n1683;
  assign n1685 = ~n594 & n1684;
  assign n1686 = ~n435 & n1685;
  assign n1687 = ~n290 & n1686;
  assign n1688 = ~n169 & ~n189;
  assign n1689 = ~n395 & n1688;
  assign n1690 = ~n601 & n1689;
  assign n1691 = ~n393 & n1690;
  assign n1692 = ~n429 & ~n518;
  assign n1693 = ~n136 & ~n299;
  assign n1694 = ~n248 & n1693;
  assign n1695 = ~n474 & n1694;
  assign n1696 = ~n155 & ~n368;
  assign n1697 = ~n363 & n1696;
  assign n1698 = n1695 & n1697;
  assign n1699 = n778 & n1698;
  assign n1700 = n1692 & n1699;
  assign n1701 = n1691 & n1700;
  assign n1702 = n1687 & n1701;
  assign n1703 = n1679 & n1702;
  assign n1704 = n1667 & n1703;
  assign n1705 = ~n168 & n1704;
  assign n1706 = ~n287 & n1705;
  assign n1707 = ~n372 & n1706;
  assign n1708 = ~n340 & n1707;
  assign n1709 = ~n466 & ~n536;
  assign n1710 = n1329 & n1709;
  assign n1711 = n1708 & n1710;
  assign n1712 = n1161 & n1711;
  assign n1713 = ~n152 & n1712;
  assign n1714 = ~n289 & n1713;
  assign n1715 = ~n146 & n1714;
  assign n1716 = ~n715 & n1715;
  assign n1717 = ~n206 & n1716;
  assign n1718 = ~n245 & n1717;
  assign n1719 = ~n158 & n1718;
  assign n1720 = ~n200 & ~n452;
  assign n1721 = ~n519 & n1720;
  assign n1722 = n1294 & n1721;
  assign n1723 = ~n123 & n1722;
  assign n1724 = ~n1246 & n1723;
  assign n1725 = ~n355 & n1724;
  assign n1726 = ~n175 & ~n228;
  assign n1727 = ~n95 & ~n666;
  assign n1728 = ~n194 & n1727;
  assign n1729 = ~n430 & n1728;
  assign n1730 = ~n274 & n1729;
  assign n1731 = ~n489 & n1730;
  assign n1732 = ~n353 & ~n1072;
  assign n1733 = ~n397 & n1732;
  assign n1734 = ~n163 & n1733;
  assign n1735 = ~n449 & n1734;
  assign n1736 = ~n490 & n1603;
  assign n1737 = ~n251 & n1736;
  assign n1738 = ~n243 & ~n637;
  assign n1739 = ~n107 & ~n883;
  assign n1740 = ~n119 & ~n495;
  assign n1741 = n1739 & n1740;
  assign n1742 = n1738 & n1741;
  assign n1743 = n1737 & n1742;
  assign n1744 = n1372 & n1743;
  assign n1745 = n1735 & n1744;
  assign n1746 = n1731 & n1745;
  assign n1747 = n1726 & n1746;
  assign n1748 = n227 & n1747;
  assign n1749 = ~n330 & n1748;
  assign n1750 = ~n426 & n1749;
  assign n1751 = ~n171 & n1750;
  assign n1752 = ~n1101 & n1751;
  assign n1753 = ~n177 & n1752;
  assign n1754 = ~n567 & n1753;
  assign n1755 = ~n233 & ~n752;
  assign n1756 = ~n144 & n1755;
  assign n1757 = ~n791 & n1756;
  assign n1758 = ~n672 & n1757;
  assign n1759 = ~n655 & n1758;
  assign n1760 = ~n232 & ~n278;
  assign n1761 = ~n424 & ~n689;
  assign n1762 = ~n469 & n1761;
  assign n1763 = ~n224 & n1762;
  assign n1764 = n1760 & n1763;
  assign n1765 = n694 & n1764;
  assign n1766 = n1759 & n1765;
  assign n1767 = n1754 & n1766;
  assign n1768 = n774 & n1767;
  assign n1769 = n1725 & n1768;
  assign n1770 = n1719 & n1769;
  assign n1771 = n1182 & n1770;
  assign n1772 = n590 & n1771;
  assign n1773 = ~n135 & n1772;
  assign n1774 = ~n400 & n1773;
  assign n1775 = ~n563 & n1774;
  assign n1776 = ~n504 & n1775;
  assign n1777 = ~n164 & n1776;
  assign n1778 = ~n325 & n1777;
  assign n1779 = ~n875 & n1778;
  assign n1780 = ~n1665 & ~n1779;
  assign n1781 = ~n655 & ~n825;
  assign n1782 = ~n189 & ~n592;
  assign n1783 = ~n154 & ~n299;
  assign n1784 = ~n1102 & n1783;
  assign n1785 = ~n163 & ~n1203;
  assign n1786 = n1784 & n1785;
  assign n1787 = n896 & n1786;
  assign n1788 = n1782 & n1787;
  assign n1789 = ~n506 & n1788;
  assign n1790 = n1755 & n1789;
  assign n1791 = ~n460 & n1790;
  assign n1792 = ~n527 & n1791;
  assign n1793 = ~n331 & n1792;
  assign n1794 = ~n689 & n1793;
  assign n1795 = ~n352 & ~n514;
  assign n1796 = ~n223 & n1795;
  assign n1797 = ~n513 & n1796;
  assign n1798 = ~n363 & n1797;
  assign n1799 = ~n335 & ~n619;
  assign n1800 = ~n438 & n1799;
  assign n1801 = n1408 & n1800;
  assign n1802 = n494 & n1801;
  assign n1803 = n1798 & n1802;
  assign n1804 = n1020 & n1803;
  assign n1805 = n515 & n1804;
  assign n1806 = n193 & n1805;
  assign n1807 = ~n136 & n1806;
  assign n1808 = ~n171 & n1807;
  assign n1809 = ~n417 & n1808;
  assign n1810 = ~n296 & n1809;
  assign n1811 = ~n274 & n1810;
  assign n1812 = ~n372 & n1811;
  assign n1813 = ~n886 & n1812;
  assign n1814 = ~n188 & n1813;
  assign n1815 = ~n469 & ~n641;
  assign n1816 = ~n203 & n1815;
  assign n1817 = ~n305 & n1816;
  assign n1818 = ~n271 & n1817;
  assign n1819 = ~n875 & n1818;
  assign n1820 = n454 & n508;
  assign n1821 = ~n563 & n1820;
  assign n1822 = ~n1104 & n1821;
  assign n1823 = ~n95 & n1822;
  assign n1824 = ~n125 & ~n158;
  assign n1825 = ~n403 & ~n602;
  assign n1826 = ~n231 & ~n504;
  assign n1827 = ~n466 & ~n777;
  assign n1828 = ~n226 & ~n1101;
  assign n1829 = n1667 & n1828;
  assign n1830 = n1827 & n1829;
  assign n1831 = n591 & n1830;
  assign n1832 = ~n1062 & n1831;
  assign n1833 = ~n290 & n1832;
  assign n1834 = ~n505 & n1833;
  assign n1835 = ~n531 & n1834;
  assign n1836 = ~n371 & n1835;
  assign n1837 = ~n569 & n1836;
  assign n1838 = ~n337 & n1837;
  assign n1839 = ~n121 & ~n536;
  assign n1840 = n962 & n1839;
  assign n1841 = ~n355 & n1840;
  assign n1842 = ~n150 & n1841;
  assign n1843 = ~n419 & n1842;
  assign n1844 = ~n603 & n1843;
  assign n1845 = n1838 & n1844;
  assign n1846 = n1826 & n1845;
  assign n1847 = n520 & n1846;
  assign n1848 = n1576 & n1847;
  assign n1849 = n826 & n1848;
  assign n1850 = n1825 & n1849;
  assign n1851 = n1824 & n1850;
  assign n1852 = ~n847 & n1851;
  assign n1853 = ~n329 & n1852;
  assign n1854 = ~n803 & n1853;
  assign n1855 = ~n571 & n1854;
  assign n1856 = ~n495 & n1855;
  assign n1857 = ~n200 & n1856;
  assign n1858 = ~n639 & n1857;
  assign n1859 = ~n492 & n1858;
  assign n1860 = ~n229 & ~n367;
  assign n1861 = ~n474 & n1860;
  assign n1862 = n1859 & n1861;
  assign n1863 = n776 & n1862;
  assign n1864 = n1823 & n1863;
  assign n1865 = n1819 & n1864;
  assign n1866 = n1814 & n1865;
  assign n1867 = n1794 & n1866;
  assign n1868 = n1531 & n1867;
  assign n1869 = n1781 & n1868;
  assign n1870 = n533 & n1869;
  assign n1871 = n282 & n1870;
  assign n1872 = n399 & n1871;
  assign n1873 = n1040 & n1872;
  assign n1874 = ~n152 & n1873;
  assign n1875 = ~n239 & n1874;
  assign n1876 = ~n287 & n1875;
  assign n1877 = ~n251 & n1876;
  assign n1878 = ~n1779 & ~n1877;
  assign n1879 = ~n165 & ~n452;
  assign n1880 = n1438 & n1879;
  assign n1881 = n1247 & n1880;
  assign n1882 = ~n398 & n1881;
  assign n1883 = ~n99 & n1882;
  assign n1884 = ~n712 & n1883;
  assign n1885 = ~n278 & ~n809;
  assign n1886 = ~n884 & n1885;
  assign n1887 = ~n245 & n1886;
  assign n1888 = ~n777 & n1887;
  assign n1889 = ~n283 & n1888;
  assign n1890 = ~n127 & n1889;
  assign n1891 = ~n136 & ~n287;
  assign n1892 = ~n298 & n1891;
  assign n1893 = ~n201 & n1892;
  assign n1894 = ~n280 & ~n667;
  assign n1895 = n618 & n1894;
  assign n1896 = ~n147 & n1895;
  assign n1897 = ~n158 & ~n511;
  assign n1898 = ~n293 & n1897;
  assign n1899 = n1896 & n1898;
  assign n1900 = n1697 & n1899;
  assign n1901 = n1345 & n1900;
  assign n1902 = n1211 & n1901;
  assign n1903 = n1039 & n1902;
  assign n1904 = n1601 & n1903;
  assign n1905 = n1476 & n1904;
  assign n1906 = n1893 & n1905;
  assign n1907 = n1890 & n1906;
  assign n1908 = n1884 & n1907;
  assign n1909 = ~n1102 & n1908;
  assign n1910 = ~n594 & n1909;
  assign n1911 = ~n419 & n1910;
  assign n1912 = ~n715 & n1911;
  assign n1913 = ~n592 & n1912;
  assign n1914 = ~n1877 & ~n1913;
  assign n1915 = ~n224 & ~n531;
  assign n1916 = ~n239 & ~n527;
  assign n1917 = ~n571 & ~n623;
  assign n1918 = ~n713 & ~n1072;
  assign n1919 = ~n329 & n1918;
  assign n1920 = ~n809 & n1919;
  assign n1921 = ~n302 & n1920;
  assign n1922 = ~n716 & n1921;
  assign n1923 = ~n132 & n1922;
  assign n1924 = ~n252 & n1923;
  assign n1925 = ~n304 & n1924;
  assign n1926 = ~n232 & ~n752;
  assign n1927 = ~n1102 & n1926;
  assign n1928 = ~n673 & n1927;
  assign n1929 = n244 & ~n426;
  assign n1930 = ~n461 & n1929;
  assign n1931 = ~n372 & n1930;
  assign n1932 = n1557 & n1931;
  assign n1933 = n874 & n1932;
  assign n1934 = n1426 & n1933;
  assign n1935 = ~n641 & n1934;
  assign n1936 = ~n514 & n1935;
  assign n1937 = ~n339 & n1936;
  assign n1938 = ~n273 & n1937;
  assign n1939 = ~n277 & n1938;
  assign n1940 = ~n325 & n1939;
  assign n1941 = ~n301 & ~n884;
  assign n1942 = ~n374 & n1941;
  assign n1943 = ~n130 & ~n299;
  assign n1944 = ~n1104 & n1943;
  assign n1945 = n989 & n1944;
  assign n1946 = n1942 & n1945;
  assign n1947 = n1940 & n1946;
  assign n1948 = n1928 & n1947;
  assign n1949 = n977 & n1948;
  assign n1950 = n538 & n1949;
  assign n1951 = ~n118 & n1950;
  assign n1952 = ~n240 & n1951;
  assign n1953 = ~n283 & n1952;
  assign n1954 = ~n791 & n1953;
  assign n1955 = ~n1203 & n1954;
  assign n1956 = ~n1010 & n1955;
  assign n1957 = ~n81 & n1956;
  assign n1958 = ~n222 & n1957;
  assign n1959 = ~n469 & ~n639;
  assign n1960 = ~n119 & n1959;
  assign n1961 = n772 & n1960;
  assign n1962 = n512 & n1961;
  assign n1963 = n1183 & n1962;
  assign n1964 = n896 & n1963;
  assign n1965 = ~n617 & n1964;
  assign n1966 = ~n367 & n1965;
  assign n1967 = ~n395 & n1966;
  assign n1968 = ~n525 & n1967;
  assign n1969 = ~n358 & n1968;
  assign n1970 = ~n121 & n221;
  assign n1971 = ~n493 & n1970;
  assign n1972 = n418 & n1248;
  assign n1973 = ~n95 & n1972;
  assign n1974 = n1971 & n1973;
  assign n1975 = n658 & n1974;
  assign n1976 = n877 & n1975;
  assign n1977 = n1969 & n1976;
  assign n1978 = n1958 & n1977;
  assign n1979 = n1925 & n1978;
  assign n1980 = n1917 & n1979;
  assign n1981 = n1916 & n1980;
  assign n1982 = n1915 & n1981;
  assign n1983 = n515 & n1982;
  assign n1984 = n1574 & n1983;
  assign n1985 = ~n558 & n1984;
  assign n1986 = ~n280 & n1985;
  assign n1987 = ~n416 & n1986;
  assign n1988 = ~n296 & n1987;
  assign n1989 = ~n505 & n1988;
  assign n1990 = ~n424 & n1989;
  assign n1991 = ~n293 & n1990;
  assign n1992 = ~n270 & n1991;
  assign n1993 = ~n1913 & ~n1992;
  assign n1994 = ~n302 & ~n1102;
  assign n1995 = ~n168 & ~n397;
  assign n1996 = ~n589 & n1995;
  assign n1997 = n1898 & n1996;
  assign n1998 = n793 & n1997;
  assign n1999 = n297 & n1998;
  assign n2000 = n1994 & n1999;
  assign n2001 = ~n1101 & n2000;
  assign n2002 = ~n205 & n2001;
  assign n2003 = ~n191 & n2002;
  assign n2004 = ~n1127 & n2003;
  assign n2005 = ~n489 & n2004;
  assign n2006 = ~n875 & n2005;
  assign n2007 = ~n492 & ~n537;
  assign n2008 = ~n667 & n2007;
  assign n2009 = ~n460 & n2008;
  assign n2010 = ~n130 & n2009;
  assign n2011 = n336 & n979;
  assign n2012 = ~n372 & n2011;
  assign n2013 = ~n340 & ~n1011;
  assign n2014 = ~n165 & ~n240;
  assign n2015 = n2013 & n2014;
  assign n2016 = n1105 & n2015;
  assign n2017 = ~n453 & n2016;
  assign n2018 = ~n355 & ~n509;
  assign n2019 = ~n147 & n2018;
  assign n2020 = ~n371 & n2019;
  assign n2021 = ~n163 & ~n716;
  assign n2022 = ~n95 & ~n746;
  assign n2023 = ~n206 & ~n364;
  assign n2024 = ~n422 & n2023;
  assign n2025 = ~n366 & n2024;
  assign n2026 = ~n222 & ~n438;
  assign n2027 = n1329 & n2026;
  assign n2028 = n529 & n2027;
  assign n2029 = n2025 & n2028;
  assign n2030 = n1691 & n2029;
  assign n2031 = n2022 & n2030;
  assign n2032 = n2021 & n2031;
  assign n2033 = n1330 & n2032;
  assign n2034 = n1668 & n2033;
  assign n2035 = n1009 & n2034;
  assign n2036 = ~n619 & n2035;
  assign n2037 = ~n192 & n2036;
  assign n2038 = ~n468 & n2037;
  assign n2039 = ~n436 & n2038;
  assign n2040 = ~n569 & n2039;
  assign n2041 = n2020 & n2040;
  assign n2042 = n2017 & n2041;
  assign n2043 = n1600 & n2042;
  assign n2044 = n2012 & n2043;
  assign n2045 = n1183 & n2044;
  assign n2046 = n2010 & n2045;
  assign n2047 = n2006 & n2046;
  assign n2048 = n720 & n2047;
  assign n2049 = ~n558 & n2048;
  assign n2050 = ~n284 & n2049;
  assign n2051 = ~n203 & n2050;
  assign n2052 = n1795 & n2051;
  assign n2053 = ~n290 & n2052;
  assign n2054 = ~n102 & n2053;
  assign n2055 = ~n424 & n2054;
  assign n2056 = ~n470 & n2055;
  assign n2057 = ~n562 & n2056;
  assign n2058 = ~n1992 & ~n2057;
  assign n2059 = ~n152 & ~n190;
  assign n2060 = n735 & n2059;
  assign n2061 = n591 & n2060;
  assign n2062 = ~n232 & n2061;
  assign n2063 = ~n809 & n2062;
  assign n2064 = ~n496 & n2063;
  assign n2065 = ~n144 & n2064;
  assign n2066 = ~n298 & n2065;
  assign n2067 = ~n337 & n2066;
  assign n2068 = ~n633 & n2067;
  assign n2069 = n1248 & n1252;
  assign n2070 = ~n289 & n2069;
  assign n2071 = ~n255 & n2070;
  assign n2072 = ~n489 & n2071;
  assign n2073 = ~n169 & ~n637;
  assign n2074 = ~n248 & n2073;
  assign n2075 = ~n1104 & n2074;
  assign n2076 = n1784 & n2075;
  assign n2077 = n812 & n2076;
  assign n2078 = n1132 & n2077;
  assign n2079 = n207 & n2078;
  assign n2080 = n1085 & n2079;
  assign n2081 = n918 & n2080;
  assign n2082 = n2072 & n2081;
  assign n2083 = n2068 & n2082;
  assign n2084 = n515 & n2083;
  assign n2085 = ~n557 & n2084;
  assign n2086 = ~n419 & n2085;
  assign n2087 = ~n396 & n2086;
  assign n2088 = ~n601 & n2087;
  assign n2089 = ~n364 & n1129;
  assign n2090 = ~n142 & ~n641;
  assign n2091 = ~n363 & ~n558;
  assign n2092 = ~n167 & ~n506;
  assign n2093 = ~n99 & ~n223;
  assign n2094 = n2092 & n2093;
  assign n2095 = n2091 & n2094;
  assign n2096 = n2090 & n2095;
  assign n2097 = n2089 & n2096;
  assign n2098 = ~n329 & n2097;
  assign n2099 = ~n150 & n2098;
  assign n2100 = ~n884 & n2099;
  assign n2101 = ~n164 & n2100;
  assign n2102 = ~n372 & n2101;
  assign n2103 = ~n393 & n2102;
  assign n2104 = ~n525 & n2103;
  assign n2105 = ~n514 & ~n713;
  assign n2106 = ~n229 & ~n667;
  assign n2107 = ~n426 & n2106;
  assign n2108 = ~n602 & n2107;
  assign n2109 = ~n115 & n2108;
  assign n2110 = ~n334 & n2109;
  assign n2111 = ~n246 & n2110;
  assign n2112 = ~n170 & n2111;
  assign n2113 = ~n226 & ~n509;
  assign n2114 = ~n1072 & n1128;
  assign n2115 = ~n146 & n2114;
  assign n2116 = n2113 & n2115;
  assign n2117 = n1643 & n2116;
  assign n2118 = n1879 & n2117;
  assign n2119 = n1012 & n2118;
  assign n2120 = n2112 & n2119;
  assign n2121 = n2021 & n2120;
  assign n2122 = n1063 & n2121;
  assign n2123 = n108 & n2122;
  assign n2124 = ~n203 & n2123;
  assign n2125 = n2105 & n2124;
  assign n2126 = ~n594 & n2125;
  assign n2127 = ~n287 & n2126;
  assign n2128 = ~n397 & ~n527;
  assign n2129 = ~n245 & n2128;
  assign n2130 = ~n567 & n2129;
  assign n2131 = ~n623 & n2130;
  assign n2132 = ~n338 & n2131;
  assign n2133 = ~n513 & ~n1062;
  assign n2134 = n475 & n2013;
  assign n2135 = n2133 & n2134;
  assign n2136 = n2132 & n2135;
  assign n2137 = n2127 & n2136;
  assign n2138 = n2104 & n2137;
  assign n2139 = n1251 & n2138;
  assign n2140 = n120 & n2139;
  assign n2141 = n2088 & n2140;
  assign n2142 = n356 & n2141;
  assign n2143 = ~n518 & n2142;
  assign n2144 = ~n151 & n2143;
  assign n2145 = ~n155 & n2144;
  assign n2146 = ~n435 & n2145;
  assign n2147 = ~n461 & n2146;
  assign n2148 = ~n326 & n2147;
  assign n2149 = ~n368 & n2148;
  assign n2150 = ~n130 & n2149;
  assign n2151 = ~n569 & n2150;
  assign n2152 = ~n655 & n2151;
  assign n2153 = ~n2057 & ~n2152;
  assign n2154 = ~n118 & ~n1072;
  assign n2155 = n1328 & n2154;
  assign n2156 = n1890 & n2155;
  assign n2157 = n1379 & n2156;
  assign n2158 = n1128 & n2157;
  assign n2159 = n2073 & n2158;
  assign n2160 = n341 & n2159;
  assign n2161 = ~n194 & n2160;
  assign n2162 = ~n1246 & n2161;
  assign n2163 = ~n803 & n2162;
  assign n2164 = ~n435 & n2163;
  assign n2165 = ~n357 & n2164;
  assign n2166 = ~n142 & n2165;
  assign n2167 = ~n271 & n2166;
  assign n2168 = ~n492 & ~n514;
  assign n2169 = ~n525 & n2168;
  assign n2170 = ~n393 & ~n980;
  assign n2171 = n356 & n2170;
  assign n2172 = ~n460 & n2171;
  assign n2173 = n156 & n1893;
  assign n2174 = ~n175 & n2173;
  assign n2175 = n747 & n773;
  assign n2176 = n1141 & n2175;
  assign n2177 = n1456 & n2176;
  assign n2178 = n2174 & n2177;
  assign n2179 = n2172 & n2178;
  assign n2180 = n757 & n2179;
  assign n2181 = n671 & n2180;
  assign n2182 = n2169 & n2181;
  assign n2183 = n1668 & n2182;
  assign n2184 = n423 & n2183;
  assign n2185 = n2167 & n2184;
  assign n2186 = n1247 & n2185;
  assign n2187 = n508 & n2186;
  assign n2188 = ~n713 & n2187;
  assign n2189 = ~n243 & n2188;
  assign n2190 = ~n2152 & ~n2189;
  assign n2191 = ~n157 & ~n276;
  assign n2192 = ~n144 & ~n1101;
  assign n2193 = n2191 & n2192;
  assign n2194 = n2154 & n2193;
  assign n2195 = n1825 & n2194;
  assign n2196 = n1550 & n2195;
  assign n2197 = n2073 & n2196;
  assign n2198 = ~n190 & n2197;
  assign n2199 = ~n278 & n2198;
  assign n2200 = ~n121 & n2199;
  assign n2201 = ~n275 & n2200;
  assign n2202 = ~n173 & n2201;
  assign n2203 = n720 & n1531;
  assign n2204 = ~n504 & n2203;
  assign n2205 = ~n271 & n2204;
  assign n2206 = ~n95 & n2205;
  assign n2207 = ~n886 & n2206;
  assign n2208 = ~n358 & n2207;
  assign n2209 = ~n714 & ~n961;
  assign n2210 = ~n147 & ~n192;
  assign n2211 = n2209 & n2210;
  assign n2212 = n887 & n2211;
  assign n2213 = ~n281 & n2212;
  assign n2214 = ~n557 & n2213;
  assign n2215 = ~n571 & n2214;
  assign n2216 = ~n228 & n2215;
  assign n2217 = ~n716 & n2216;
  assign n2218 = ~n194 & ~n619;
  assign n2219 = ~n825 & n2218;
  assign n2220 = ~n273 & ~n506;
  assign n2221 = n595 & n2220;
  assign n2222 = n2093 & n2221;
  assign n2223 = n1069 & n2222;
  assign n2224 = ~n354 & n2223;
  assign n2225 = ~n803 & n2224;
  assign n2226 = ~n367 & n2225;
  assign n2227 = ~n146 & n2226;
  assign n2228 = ~n286 & n2227;
  assign n2229 = ~n245 & n2228;
  assign n2230 = ~n236 & ~n460;
  assign n2231 = n133 & n2230;
  assign n2232 = n1942 & n2231;
  assign n2233 = ~n752 & n2232;
  assign n2234 = ~n189 & n2233;
  assign n2235 = ~n417 & n2234;
  assign n2236 = ~n453 & n2235;
  assign n2237 = ~n394 & n2236;
  assign n2238 = ~n352 & ~n420;
  assign n2239 = ~n505 & n2238;
  assign n2240 = ~n163 & n2239;
  assign n2241 = ~n107 & ~n563;
  assign n2242 = n1763 & n2241;
  assign n2243 = n2240 & n2242;
  assign n2244 = n2237 & n2243;
  assign n2245 = n808 & n2244;
  assign n2246 = n2229 & n2245;
  assign n2247 = n1994 & n2246;
  assign n2248 = n2219 & n2247;
  assign n2249 = n116 & n2248;
  assign n2250 = n1389 & n2249;
  assign n2251 = ~n136 & n2250;
  assign n2252 = ~n713 & n2251;
  assign n2253 = ~n641 & n2252;
  assign n2254 = ~n292 & n2253;
  assign n2255 = ~n396 & n2254;
  assign n2256 = ~n248 & n2255;
  assign n2257 = ~n290 & n2256;
  assign n2258 = ~n567 & n2257;
  assign n2259 = n618 & n1827;
  assign n2260 = ~n239 & n2259;
  assign n2261 = ~n513 & n2260;
  assign n2262 = ~n429 & n2261;
  assign n2263 = ~n746 & ~n809;
  assign n2264 = ~n161 & n202;
  assign n2265 = ~n672 & n2264;
  assign n2266 = n526 & n732;
  assign n2267 = ~n237 & n2266;
  assign n2268 = n2265 & n2267;
  assign n2269 = n535 & n2268;
  assign n2270 = n1155 & n2269;
  assign n2271 = ~n623 & n2270;
  assign n2272 = ~n712 & n2271;
  assign n2273 = ~n436 & n2272;
  assign n2274 = ~n225 & n2273;
  assign n2275 = ~n158 & n2274;
  assign n2276 = ~n496 & ~n601;
  assign n2277 = ~n152 & n2276;
  assign n2278 = ~n357 & n2277;
  assign n2279 = n2275 & n2278;
  assign n2280 = n365 & n2279;
  assign n2281 = n2263 & n2280;
  assign n2282 = n2262 & n2281;
  assign n2283 = n1268 & n2282;
  assign n2284 = n2258 & n2283;
  assign n2285 = n2217 & n2284;
  assign n2286 = n2208 & n2285;
  assign n2287 = n2202 & n2286;
  assign n2288 = n510 & n2287;
  assign n2289 = ~n355 & n2288;
  assign n2290 = ~n255 & n2289;
  assign n2291 = ~n620 & n2290;
  assign n2292 = ~n2189 & ~n2291;
  assign n2293 = ~n243 & ~n367;
  assign n2294 = ~n228 & n2293;
  assign n2295 = ~n537 & n2294;
  assign n2296 = ~n470 & n2295;
  assign n2297 = ~n146 & ~n460;
  assign n2298 = n827 & n2297;
  assign n2299 = ~n847 & n2298;
  assign n2300 = ~n150 & n2299;
  assign n2301 = ~n290 & n2300;
  assign n2302 = n1131 & n1476;
  assign n2303 = ~n746 & n2302;
  assign n2304 = n1025 & n2303;
  assign n2305 = n1533 & n2304;
  assign n2306 = n816 & n2305;
  assign n2307 = n207 & n2306;
  assign n2308 = n2091 & n2307;
  assign n2309 = n2301 & n2308;
  assign n2310 = n2296 & n2309;
  assign n2311 = n2169 & n2310;
  assign n2312 = n1825 & n2311;
  assign n2313 = ~n229 & n2312;
  assign n2314 = ~n777 & n2313;
  assign n2315 = ~n287 & n2314;
  assign n2316 = ~n603 & n2315;
  assign n2317 = ~n1104 & n2316;
  assign n2318 = ~n171 & ~n354;
  assign n2319 = ~n280 & n2318;
  assign n2320 = ~n275 & n2319;
  assign n2321 = ~n292 & n2320;
  assign n2322 = ~n416 & n2321;
  assign n2323 = ~n192 & n2322;
  assign n2324 = ~n164 & n2323;
  assign n2325 = ~n567 & n2324;
  assign n2326 = ~n301 & n437;
  assign n2327 = ~n339 & n2326;
  assign n2328 = ~n357 & n2327;
  assign n2329 = ~n657 & n2328;
  assign n2330 = ~n188 & n2329;
  assign n2331 = ~n601 & ~n667;
  assign n2332 = ~n337 & n2331;
  assign n2333 = ~n167 & ~n331;
  assign n2334 = ~n252 & n2333;
  assign n2335 = n887 & n2334;
  assign n2336 = n2332 & n2335;
  assign n2337 = n632 & n2336;
  assign n2338 = n2330 & n2337;
  assign n2339 = n238 & n2338;
  assign n2340 = n2325 & n2339;
  assign n2341 = n896 & n2340;
  assign n2342 = ~n420 & n2341;
  assign n2343 = ~n353 & n2342;
  assign n2344 = ~n155 & n2343;
  assign n2345 = ~n1127 & n2344;
  assign n2346 = ~n563 & ~n673;
  assign n2347 = ~n175 & n2346;
  assign n2348 = ~n468 & ~n961;
  assign n2349 = ~n589 & ~n1246;
  assign n2350 = n1636 & n1739;
  assign n2351 = n2349 & n2350;
  assign n2352 = n2348 & n2351;
  assign n2353 = n241 & n2352;
  assign n2354 = ~n1102 & n2353;
  assign n2355 = n2347 & n2354;
  assign n2356 = ~n327 & n2355;
  assign n2357 = ~n594 & n2356;
  assign n2358 = ~n430 & n2357;
  assign n2359 = ~n1203 & n2358;
  assign n2360 = ~n474 & n2359;
  assign n2361 = ~n302 & ~n532;
  assign n2362 = ~n91 & ~n518;
  assign n2363 = ~n142 & n2362;
  assign n2364 = n2361 & n2363;
  assign n2365 = ~n281 & n2364;
  assign n2366 = ~n147 & n2365;
  assign n2367 = ~n791 & n2366;
  assign n2368 = ~n493 & n2367;
  assign n2369 = ~n358 & n2368;
  assign n2370 = ~n875 & n2369;
  assign n2371 = ~n328 & ~n569;
  assign n2372 = n793 & n1839;
  assign n2373 = n308 & n2372;
  assign n2374 = n2371 & n2373;
  assign n2375 = n2370 & n2374;
  assign n2376 = n2360 & n2375;
  assign n2377 = n2345 & n2376;
  assign n2378 = n2317 & n2377;
  assign n2379 = n1667 & n2378;
  assign n2380 = n937 & n2379;
  assign n2381 = n1252 & n2380;
  assign n2382 = ~n462 & n2381;
  assign n2383 = n1021 & n2382;
  assign n2384 = ~n715 & n2383;
  assign n2385 = ~n157 & n2384;
  assign n2386 = ~n325 & n2385;
  assign n2387 = ~n886 & n2386;
  assign n2388 = ~n231 & n2387;
  assign n2389 = ~n2291 & ~n2388;
  assign n2390 = ~n173 & ~n564;
  assign n2391 = n362 & n2390;
  assign n2392 = n1879 & n2391;
  assign n2393 = n1380 & n2392;
  assign n2394 = n1761 & n2393;
  assign n2395 = ~n123 & n2394;
  assign n2396 = n1108 & n2395;
  assign n2397 = ~n511 & n2396;
  assign n2398 = ~n118 & n2397;
  assign n2399 = ~n417 & n2398;
  assign n2400 = ~n290 & n2399;
  assign n2401 = ~n777 & n2400;
  assign n2402 = ~n537 & n2401;
  assign n2403 = ~n200 & n2402;
  assign n2404 = ~n272 & n2403;
  assign n2405 = ~n1127 & n2404;
  assign n2406 = ~n99 & ~n451;
  assign n2407 = ~n273 & ~n292;
  assign n2408 = ~n883 & n2407;
  assign n2409 = ~n428 & n2408;
  assign n2410 = ~n147 & ~n271;
  assign n2411 = n1324 & n2410;
  assign n2412 = ~n639 & n2411;
  assign n2413 = ~n825 & n2412;
  assign n2414 = ~n145 & n2413;
  assign n2415 = ~n240 & n2414;
  assign n2416 = ~n372 & n2415;
  assign n2417 = ~n589 & n2416;
  assign n2418 = ~n637 & ~n1102;
  assign n2419 = ~n205 & n2418;
  assign n2420 = ~n1203 & n2419;
  assign n2421 = ~n470 & n2420;
  assign n2422 = ~n592 & n2421;
  assign n2423 = ~n119 & ~n142;
  assign n2424 = ~n223 & ~n419;
  assign n2425 = ~n248 & ~n1062;
  assign n2426 = ~n368 & n2425;
  assign n2427 = n156 & ~n932;
  assign n2428 = n2426 & n2427;
  assign n2429 = n2424 & n2428;
  assign n2430 = n2423 & n2429;
  assign n2431 = n2422 & n2430;
  assign n2432 = n1131 & n2431;
  assign n2433 = n2417 & n2432;
  assign n2434 = n1247 & n2433;
  assign n2435 = ~n236 & n2434;
  assign n2436 = ~n242 & n2435;
  assign n2437 = ~n284 & n2436;
  assign n2438 = ~n130 & n2437;
  assign n2439 = ~n449 & n2438;
  assign n2440 = n288 & n2439;
  assign n2441 = ~n429 & n2440;
  assign n2442 = ~n301 & ~n712;
  assign n2443 = ~n791 & n2442;
  assign n2444 = ~n425 & n2443;
  assign n2445 = ~n657 & n2444;
  assign n2446 = n2441 & n2445;
  assign n2447 = n2409 & n2446;
  assign n2448 = n790 & n2447;
  assign n2449 = n2040 & n2448;
  assign n2450 = n665 & n2449;
  assign n2451 = n604 & n2450;
  assign n2452 = n2406 & n2451;
  assign n2453 = n1667 & n2452;
  assign n2454 = n399 & n2453;
  assign n2455 = n2068 & n2454;
  assign n2456 = n2405 & n2455;
  assign n2457 = ~n713 & n2456;
  assign n2458 = ~n233 & n2457;
  assign n2459 = ~n461 & n2458;
  assign n2460 = ~n157 & n2459;
  assign n2461 = ~n623 & n2460;
  assign n2462 = ~n338 & n2461;
  assign n2463 = ~n532 & n2462;
  assign n2464 = ~n666 & n2463;
  assign n2465 = ~n2388 & ~n2464;
  assign n2466 = ~n255 & ~n617;
  assign n2467 = ~n305 & ~n451;
  assign n2468 = ~n366 & ~n689;
  assign n2469 = n202 & ~n495;
  assign n2470 = ~n252 & n2469;
  assign n2471 = n990 & n2470;
  assign n2472 = n899 & n2471;
  assign n2473 = n2468 & n2472;
  assign n2474 = n2348 & n2473;
  assign n2475 = n2467 & n2474;
  assign n2476 = n193 & n2475;
  assign n2477 = n2466 & n2476;
  assign n2478 = ~n396 & n2477;
  assign n2479 = ~n290 & n2478;
  assign n2480 = ~n283 & n2479;
  assign n2481 = ~n525 & n2480;
  assign n2482 = ~n158 & n2481;
  assign n2483 = ~n655 & n2482;
  assign n2484 = ~n167 & ~n430;
  assign n2485 = ~n490 & ~n514;
  assign n2486 = ~n374 & n2485;
  assign n2487 = ~n603 & n2486;
  assign n2488 = n365 & n1204;
  assign n2489 = n300 & n2488;
  assign n2490 = n2487 & n2489;
  assign n2491 = n1915 & n2490;
  assign n2492 = n621 & n2491;
  assign n2493 = n896 & n2492;
  assign n2494 = n885 & n2493;
  assign n2495 = ~n1072 & n2494;
  assign n2496 = ~n111 & n2495;
  assign n2497 = ~n809 & n2496;
  assign n2498 = ~n121 & n2497;
  assign n2499 = ~n1010 & n2498;
  assign n2500 = ~n771 & n2499;
  assign n2501 = ~n460 & ~n594;
  assign n2502 = ~n206 & n2501;
  assign n2503 = ~n243 & n2502;
  assign n2504 = ~n657 & n2503;
  assign n2505 = ~n161 & n2504;
  assign n2506 = ~n672 & n2505;
  assign n2507 = ~n163 & ~n1246;
  assign n2508 = ~n420 & ~n504;
  assign n2509 = n642 & n2508;
  assign n2510 = ~n435 & n2509;
  assign n2511 = ~n292 & n2510;
  assign n2512 = ~n519 & n2511;
  assign n2513 = ~n232 & n282;
  assign n2514 = ~n713 & n2513;
  assign n2515 = ~n231 & n2514;
  assign n2516 = n351 & n2515;
  assign n2517 = n2512 & n2516;
  assign n2518 = n2507 & n2517;
  assign n2519 = n2439 & n2518;
  assign n2520 = n2506 & n2519;
  assign n2521 = n2500 & n2520;
  assign n2522 = n2484 & n2521;
  assign n2523 = n720 & n2522;
  assign n2524 = n2483 & n2523;
  assign n2525 = ~n189 & n2524;
  assign n2526 = ~n239 & n2525;
  assign n2527 = ~n417 & n2526;
  assign n2528 = ~n226 & n2527;
  assign n2529 = ~n438 & n2528;
  assign n2530 = ~n563 & n2529;
  assign n2531 = ~n791 & n2530;
  assign n2532 = ~n295 & n2531;
  assign n2533 = ~n293 & n2532;
  assign n2534 = ~n2464 & ~n2533;
  assign n2535 = ~n248 & ~n327;
  assign n2536 = ~n91 & n2535;
  assign n2537 = ~n273 & n2536;
  assign n2538 = n624 & n2537;
  assign n2539 = ~n961 & n2538;
  assign n2540 = ~n130 & n2539;
  assign n2541 = ~n225 & n2540;
  assign n2542 = ~n252 & n2541;
  assign n2543 = ~n95 & n2542;
  assign n2544 = ~n398 & ~n594;
  assign n2545 = ~n242 & ~n505;
  assign n2546 = ~n157 & n2545;
  assign n2547 = n2427 & n2546;
  assign n2548 = n2544 & n2547;
  assign n2549 = n2170 & n2548;
  assign n2550 = ~n255 & n2549;
  assign n2551 = ~n619 & n2550;
  assign n2552 = ~n287 & n2551;
  assign n2553 = ~n306 & n2552;
  assign n2554 = ~n371 & n2553;
  assign n2555 = ~n231 & n2554;
  assign n2556 = ~n239 & ~n633;
  assign n2557 = n638 & n2556;
  assign n2558 = n989 & n2557;
  assign n2559 = n1879 & n2558;
  assign n2560 = n844 & n2559;
  assign n2561 = n1202 & n2560;
  assign n2562 = n2555 & n2561;
  assign n2563 = n2543 & n2562;
  assign n2564 = n1379 & n2563;
  assign n2565 = n1389 & n2564;
  assign n2566 = ~n397 & n2565;
  assign n2567 = ~n752 & n2566;
  assign n2568 = ~n334 & n2567;
  assign n2569 = ~n107 & n2568;
  assign n2570 = ~n716 & n2569;
  assign n2571 = ~n569 & n2570;
  assign n2572 = ~n2533 & ~n2571;
  assign n2573 = ~n325 & ~n883;
  assign n2574 = ~n427 & ~n617;
  assign n2575 = ~n254 & n2574;
  assign n2576 = ~n803 & n2575;
  assign n2577 = ~n228 & n2576;
  assign n2578 = ~n191 & n2577;
  assign n2579 = ~n283 & n2578;
  assign n2580 = ~n366 & n2579;
  assign n2581 = ~n489 & n2580;
  assign n2582 = ~n363 & ~n875;
  assign n2583 = ~n509 & ~n623;
  assign n2584 = ~n398 & ~n468;
  assign n2585 = n2090 & n2584;
  assign n2586 = ~n847 & n2585;
  assign n2587 = ~n175 & n2586;
  assign n2588 = ~n223 & n2587;
  assign n2589 = ~n568 & n2588;
  assign n2590 = ~n340 & n2589;
  assign n2591 = ~n1127 & n2590;
  assign n2592 = ~n240 & ~n245;
  assign n2593 = ~n1203 & n2592;
  assign n2594 = n873 & n1180;
  assign n2595 = ~n95 & n2594;
  assign n2596 = n2593 & n2595;
  assign n2597 = n2349 & n2596;
  assign n2598 = n1839 & n2597;
  assign n2599 = n977 & n2598;
  assign n2600 = ~n115 & n2599;
  assign n2601 = ~n514 & n2600;
  assign n2602 = ~n435 & n2601;
  assign n2603 = ~n225 & n2602;
  assign n2604 = ~n532 & n2603;
  assign n2605 = ~n81 & n2604;
  assign n2606 = ~n169 & ~n537;
  assign n2607 = ~n525 & n2606;
  assign n2608 = ~n461 & ~n504;
  assign n2609 = n1800 & n2608;
  assign n2610 = n2607 & n2609;
  assign n2611 = n595 & n2610;
  assign n2612 = n790 & n2611;
  assign n2613 = n2605 & n2612;
  assign n2614 = n2591 & n2613;
  assign n2615 = n1602 & n2614;
  assign n2616 = n2583 & n2615;
  assign n2617 = n2582 & n2616;
  assign n2618 = ~n364 & n2617;
  assign n2619 = ~n168 & n2618;
  assign n2620 = ~n352 & n2619;
  assign n2621 = ~n118 & n2620;
  assign n2622 = ~n424 & n2621;
  assign n2623 = ~n673 & n2622;
  assign n2624 = ~n511 & n616;
  assign n2625 = ~n130 & n2624;
  assign n2626 = ~n194 & ~n558;
  assign n2627 = ~n714 & n2626;
  assign n2628 = n2625 & n2627;
  assign n2629 = n2371 & n2628;
  assign n2630 = ~n242 & n2629;
  assign n2631 = ~n357 & n2630;
  assign n2632 = ~n712 & n2631;
  assign n2633 = ~n123 & ~n393;
  assign n2634 = ~n177 & ~n201;
  assign n2635 = ~n252 & n2634;
  assign n2636 = ~n206 & n2635;
  assign n2637 = ~n358 & n2636;
  assign n2638 = n1578 & n1828;
  assign n2639 = n2637 & n2638;
  assign n2640 = n1738 & n2639;
  assign n2641 = n1419 & n2640;
  assign n2642 = n811 & n2641;
  assign n2643 = n2633 & n2642;
  assign n2644 = n933 & n2643;
  assign n2645 = n2484 & n2644;
  assign n2646 = ~n397 & n2645;
  assign n2647 = ~n102 & n2646;
  assign n2648 = ~n237 & n2647;
  assign n2649 = ~n562 & n2648;
  assign n2650 = ~n655 & n2649;
  assign n2651 = ~n91 & ~n505;
  assign n2652 = n282 & n2651;
  assign n2653 = ~n527 & n2652;
  assign n2654 = ~n420 & ~n602;
  assign n2655 = ~n173 & n2654;
  assign n2656 = ~n493 & n2655;
  assign n2657 = n2653 & n2656;
  assign n2658 = n2650 & n2657;
  assign n2659 = n2632 & n2658;
  assign n2660 = n2623 & n2659;
  assign n2661 = n2581 & n2660;
  assign n2662 = n2573 & n2661;
  assign n2663 = n159 & n2662;
  assign n2664 = n979 & n2663;
  assign n2665 = n720 & n2664;
  assign n2666 = ~n1072 & n2665;
  assign n2667 = ~n469 & n2666;
  assign n2668 = ~n518 & n2667;
  assign n2669 = ~n980 & n2668;
  assign n2670 = ~n277 & n2669;
  assign n2671 = ~n564 & n2670;
  assign n2672 = ~n371 & n2671;
  assign n2673 = ~n188 & n2672;
  assign n2674 = ~n231 & n2673;
  assign n2675 = ~n2571 & ~n2674;
  assign n2676 = ~n355 & ~n504;
  assign n2677 = ~n240 & n2676;
  assign n2678 = ~n304 & n2677;
  assign n2679 = n128 & n1121;
  assign n2680 = ~n603 & n2679;
  assign n2681 = ~n1203 & n2680;
  assign n2682 = ~n531 & n2681;
  assign n2683 = ~n222 & ~n287;
  assign n2684 = ~n115 & n2683;
  assign n2685 = n2390 & n2684;
  assign n2686 = n2133 & n2685;
  assign n2687 = n1387 & n2686;
  assign n2688 = n2682 & n2687;
  assign n2689 = n2325 & n2688;
  assign n2690 = n1182 & n2689;
  assign n2691 = n979 & n2690;
  assign n2692 = n2583 & n2691;
  assign n2693 = ~n169 & n2692;
  assign n2694 = ~n396 & n2693;
  assign n2695 = ~n1104 & n2694;
  assign n2696 = ~n883 & n2695;
  assign n2697 = ~n95 & n2696;
  assign n2698 = ~n422 & ~n525;
  assign n2699 = ~n571 & ~n809;
  assign n2700 = ~n514 & n2699;
  assign n2701 = ~n339 & n2700;
  assign n2702 = ~n233 & n2701;
  assign n2703 = ~n248 & n2702;
  assign n2704 = ~n601 & ~n875;
  assign n2705 = ~n175 & ~n295;
  assign n2706 = n1636 & n2705;
  assign n2707 = n2704 & n2706;
  assign n2708 = n2507 & n2707;
  assign n2709 = ~n1011 & n2708;
  assign n2710 = ~n495 & n2709;
  assign n2711 = ~n118 & n2710;
  assign n2712 = ~n400 & n2711;
  assign n2713 = ~n777 & n2712;
  assign n2714 = ~n394 & n2713;
  assign n2715 = ~n886 & n2714;
  assign n2716 = ~n270 & n2715;
  assign n2717 = ~n453 & n1782;
  assign n2718 = ~n306 & n2717;
  assign n2719 = ~n249 & n2718;
  assign n2720 = ~n255 & ~n563;
  assign n2721 = ~n86 & n2720;
  assign n2722 = n2303 & n2721;
  assign n2723 = n2230 & n2722;
  assign n2724 = n2719 & n2723;
  assign n2725 = n2650 & n2724;
  assign n2726 = n2716 & n2725;
  assign n2727 = n2703 & n2726;
  assign n2728 = n2698 & n2727;
  assign n2729 = n1183 & n2728;
  assign n2730 = n2697 & n2729;
  assign n2731 = n2678 & n2730;
  assign n2732 = n937 & n2731;
  assign n2733 = ~n619 & n2732;
  assign n2734 = ~n639 & n2733;
  assign n2735 = ~n200 & n2734;
  assign n2736 = ~n1010 & n2735;
  assign n2737 = ~n2674 & ~n2736;
  assign n2738 = ~n229 & ~n1246;
  assign n2739 = ~n334 & ~n656;
  assign n2740 = ~n151 & ~n171;
  assign n2741 = ~n355 & n804;
  assign n2742 = ~n875 & n2741;
  assign n2743 = n2740 & n2742;
  assign n2744 = n2739 & n2743;
  assign n2745 = n1128 & n2744;
  assign n2746 = ~n135 & n2745;
  assign n2747 = ~n809 & n2746;
  assign n2748 = ~n223 & n2747;
  assign n2749 = ~n715 & n2748;
  assign n2750 = ~n438 & n2749;
  assign n2751 = ~n252 & n2750;
  assign n2752 = ~n436 & ~n567;
  assign n2753 = ~n400 & n520;
  assign n2754 = n2752 & n2753;
  assign n2755 = n2445 & n2754;
  assign n2756 = n2544 & n2755;
  assign n2757 = n494 & n2756;
  assign n2758 = ~n152 & ~n617;
  assign n2759 = ~n118 & n2758;
  assign n2760 = n1314 & n2759;
  assign n2761 = n2757 & n2760;
  assign n2762 = n2751 & n2761;
  assign n2763 = n2738 & n2762;
  assign n2764 = n1253 & n2763;
  assign n2765 = n2651 & n2764;
  assign n2766 = n507 & n2765;
  assign n2767 = ~n254 & n2766;
  assign n2768 = ~n328 & n2767;
  assign n2769 = ~n299 & n2768;
  assign n2770 = ~n568 & n2769;
  assign n2771 = ~n243 & n2770;
  assign n2772 = ~n531 & n2771;
  assign n2773 = ~n746 & ~n1011;
  assign n2774 = ~n402 & n2773;
  assign n2775 = ~n305 & n2774;
  assign n2776 = ~n825 & n2775;
  assign n2777 = ~n672 & n2776;
  assign n2778 = ~n371 & n2777;
  assign n2779 = n566 & n1727;
  assign n2780 = ~n426 & n2779;
  assign n2781 = ~n367 & n2780;
  assign n2782 = ~n145 & n2781;
  assign n2783 = n418 & ~n492;
  assign n2784 = ~n245 & n2783;
  assign n2785 = n632 & n2784;
  assign n2786 = n204 & n2785;
  assign n2787 = n2782 & n2786;
  assign n2788 = n2778 & n2787;
  assign n2789 = n1994 & n2788;
  assign n2790 = n515 & n2789;
  assign n2791 = n1237 & n2790;
  assign n2792 = n634 & n2791;
  assign n2793 = ~n416 & n2792;
  assign n2794 = ~n714 & n2793;
  assign n2795 = ~n393 & n2794;
  assign n2796 = ~n489 & n2795;
  assign n2797 = n1025 & n1602;
  assign n2798 = n1426 & n2797;
  assign n2799 = n654 & n2798;
  assign n2800 = ~n1072 & n2799;
  assign n2801 = ~n509 & n2800;
  assign n2802 = ~n147 & n2801;
  assign n2803 = ~n130 & n2802;
  assign n2804 = ~n525 & n2803;
  assign n2805 = ~n127 & n2804;
  assign n2806 = ~n655 & n2805;
  assign n2807 = ~n132 & ~n325;
  assign n2808 = ~n194 & ~n886;
  assign n2809 = ~n293 & ~n372;
  assign n2810 = ~n164 & n2073;
  assign n2811 = ~n277 & n2810;
  assign n2812 = n1828 & n2811;
  assign n2813 = n2809 & n2812;
  assign n2814 = n2808 & n2813;
  assign n2815 = n2807 & n2814;
  assign n2816 = n1709 & n2815;
  assign n2817 = n2806 & n2816;
  assign n2818 = n2796 & n2817;
  assign n2819 = n2772 & n2818;
  assign n2820 = n789 & n2819;
  assign n2821 = n1577 & n2820;
  assign n2822 = n1917 & n2821;
  assign n2823 = n533 & n2822;
  assign n2824 = n421 & n2823;
  assign n2825 = n2276 & n2824;
  assign n2826 = ~n284 & n2825;
  assign n2827 = ~n146 & n2826;
  assign n2828 = ~n331 & n2827;
  assign n2829 = ~n274 & n2828;
  assign n2830 = n2674 & ~n2736;
  assign n2831 = ~n2829 & n2830;
  assign n2832 = ~n2737 & ~n2831;
  assign n2833 = n2571 & n2674;
  assign n2834 = ~n2675 & ~n2833;
  assign n2835 = ~n2832 & n2834;
  assign n2836 = ~n2675 & ~n2835;
  assign n2837 = n2533 & n2571;
  assign n2838 = ~n2572 & ~n2837;
  assign n2839 = ~n2836 & n2838;
  assign n2840 = ~n2572 & ~n2839;
  assign n2841 = n2464 & n2533;
  assign n2842 = ~n2534 & ~n2841;
  assign n2843 = ~n2840 & n2842;
  assign n2844 = ~n2534 & ~n2843;
  assign n2845 = n2388 & n2464;
  assign n2846 = ~n2465 & ~n2845;
  assign n2847 = ~n2844 & n2846;
  assign n2848 = ~n2465 & ~n2847;
  assign n2849 = n2291 & n2388;
  assign n2850 = ~n2389 & ~n2849;
  assign n2851 = ~n2848 & n2850;
  assign n2852 = ~n2389 & ~n2851;
  assign n2853 = n2189 & n2291;
  assign n2854 = ~n2292 & ~n2853;
  assign n2855 = ~n2852 & n2854;
  assign n2856 = ~n2292 & ~n2855;
  assign n2857 = n2152 & n2189;
  assign n2858 = ~n2190 & ~n2857;
  assign n2859 = ~n2856 & n2858;
  assign n2860 = ~n2190 & ~n2859;
  assign n2861 = n2057 & n2152;
  assign n2862 = ~n2153 & ~n2861;
  assign n2863 = ~n2860 & n2862;
  assign n2864 = ~n2153 & ~n2863;
  assign n2865 = n1992 & n2057;
  assign n2866 = ~n2058 & ~n2865;
  assign n2867 = ~n2864 & n2866;
  assign n2868 = ~n2058 & ~n2867;
  assign n2869 = n1913 & n1992;
  assign n2870 = ~n1993 & ~n2869;
  assign n2871 = ~n2868 & n2870;
  assign n2872 = ~n1993 & ~n2871;
  assign n2873 = n1877 & n1913;
  assign n2874 = ~n1914 & ~n2873;
  assign n2875 = ~n2872 & n2874;
  assign n2876 = ~n1914 & ~n2875;
  assign n2877 = n1779 & n1877;
  assign n2878 = ~n1878 & ~n2877;
  assign n2879 = ~n2876 & n2878;
  assign n2880 = ~n1878 & ~n2879;
  assign n2881 = n1665 & n1779;
  assign n2882 = ~n1780 & ~n2881;
  assign n2883 = ~n2880 & n2882;
  assign n2884 = ~n1780 & ~n2883;
  assign n2885 = n1572 & n1665;
  assign n2886 = ~n1666 & ~n2885;
  assign n2887 = ~n2884 & n2886;
  assign n2888 = ~n1666 & ~n2887;
  assign n2889 = n1472 & n1572;
  assign n2890 = ~n1573 & ~n2889;
  assign n2891 = ~n2888 & n2890;
  assign n2892 = ~n1573 & ~n2891;
  assign n2893 = n1364 & n1472;
  assign n2894 = ~n1473 & ~n2893;
  assign n2895 = ~n2892 & n2894;
  assign n2896 = ~n1473 & ~n2895;
  assign n2897 = n1235 & n1364;
  assign n2898 = ~n1365 & ~n2897;
  assign n2899 = ~n2896 & n2898;
  assign n2900 = ~n1365 & ~n2899;
  assign n2901 = n1178 & n1235;
  assign n2902 = ~n1236 & ~n2901;
  assign n2903 = ~n2900 & n2902;
  assign n2904 = ~n1236 & ~n2903;
  assign n2905 = n1060 & n1178;
  assign n2906 = ~n1179 & ~n2905;
  assign n2907 = ~n2904 & n2906;
  assign n2908 = ~n1179 & ~n2907;
  assign n2909 = n958 & n1060;
  assign n2910 = ~n1061 & ~n2909;
  assign n2911 = ~n2908 & n2910;
  assign n2912 = ~n1061 & ~n2911;
  assign n2913 = n867 & n958;
  assign n2914 = ~n959 & ~n2913;
  assign n2915 = ~n2912 & n2914;
  assign n2916 = ~n959 & ~n2915;
  assign n2917 = n710 & n867;
  assign n2918 = ~n868 & ~n2917;
  assign n2919 = ~n2916 & n2918;
  assign n2920 = ~n868 & ~n2919;
  assign n2921 = n587 & n710;
  assign n2922 = ~n711 & ~n2921;
  assign n2923 = ~n2920 & n2922;
  assign n2924 = ~n711 & ~n2923;
  assign n2925 = n392 & n587;
  assign n2926 = ~n588 & ~n2925;
  assign n2927 = ~n2924 & n2926;
  assign n2928 = ~n588 & ~n2927;
  assign n2929 = ~n206 & ~n327;
  assign n2930 = ~n468 & n2929;
  assign n2931 = ~n655 & n2930;
  assign n2932 = n2090 & n2931;
  assign n2933 = ~n1072 & n2932;
  assign n2934 = ~n557 & n2933;
  assign n2935 = ~n426 & n2934;
  assign n2936 = ~n637 & n2935;
  assign n2937 = ~n306 & n2936;
  assign n2938 = ~n672 & n2937;
  assign n2939 = ~n337 & n2938;
  assign n2940 = ~n771 & n2939;
  assign n2941 = ~n149 & n1556;
  assign n2942 = ~n568 & n2941;
  assign n2943 = ~n99 & n2942;
  assign n2944 = n990 & n1408;
  assign n2945 = n2943 & n2944;
  assign n2946 = n2940 & n2945;
  assign n2947 = n2219 & n2946;
  assign n2948 = n1180 & n2947;
  assign n2949 = ~n301 & n2948;
  assign n2950 = ~n276 & n2949;
  assign n2951 = ~n355 & n2950;
  assign n2952 = ~n335 & n2951;
  assign n2953 = ~n639 & n2952;
  assign n2954 = ~n714 & n2953;
  assign n2955 = ~n274 & n2954;
  assign n2956 = ~n240 & n2955;
  assign n2957 = ~n277 & n2956;
  assign n2958 = ~n325 & n2957;
  assign n2959 = n2263 & n2752;
  assign n2960 = ~n462 & n2959;
  assign n2961 = ~n980 & n2960;
  assign n2962 = ~n713 & n1760;
  assign n2963 = ~n281 & n2962;
  assign n2964 = n832 & n1423;
  assign n2965 = n2230 & n2964;
  assign n2966 = n2963 & n2965;
  assign n2967 = n2961 & n2966;
  assign n2968 = n1916 & n2967;
  assign n2969 = n2021 & n2968;
  assign n2970 = n288 & n2969;
  assign n2971 = n533 & n2970;
  assign n2972 = n1825 & n2971;
  assign n2973 = n2466 & n2972;
  assign n2974 = ~n594 & n2973;
  assign n2975 = ~n470 & n2974;
  assign n2976 = ~n592 & n2975;
  assign n2977 = ~n666 & n2976;
  assign n2978 = ~n489 & n2977;
  assign n2979 = ~n249 & n2978;
  assign n2980 = ~n171 & n2409;
  assign n2981 = ~n305 & n2980;
  assign n2982 = ~n102 & n2981;
  assign n2983 = ~n331 & n2982;
  assign n2984 = ~n283 & n2983;
  assign n2985 = ~n372 & n2984;
  assign n2986 = ~n1010 & n2985;
  assign n2987 = ~n519 & n2986;
  assign n2988 = n634 & n1009;
  assign n2989 = ~n289 & n2988;
  assign n2990 = ~n531 & n2989;
  assign n2991 = ~n352 & n421;
  assign n2992 = ~n338 & n2991;
  assign n2993 = ~n121 & ~n177;
  assign n2994 = ~n398 & n2993;
  assign n2995 = ~n115 & n2994;
  assign n2996 = n2113 & n2995;
  assign n2997 = n2992 & n2996;
  assign n2998 = n2990 & n2997;
  assign n2999 = n1823 & n2998;
  assign n3000 = n2987 & n2999;
  assign n3001 = n2979 & n3000;
  assign n3002 = n244 & n3001;
  assign n3003 = n2958 & n3002;
  assign n3004 = n590 & n3003;
  assign n3005 = n1389 & n3004;
  assign n3006 = ~n136 & n3005;
  assign n3007 = ~n506 & n3006;
  assign n3008 = ~n357 & n3007;
  assign n3009 = ~n326 & n3008;
  assign n3010 = ~n1203 & n3009;
  assign n3011 = ~n200 & n3010;
  assign n3012 = ~n371 & n3011;
  assign n3013 = ~n392 & ~n3012;
  assign n3014 = n392 & n3012;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = ~n2928 & n3015;
  assign n3017 = n2928 & ~n3015;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = n75 & n3018;
  assign n3020 = ~ a[31]  & ~n74;
  assign n3021 = ~n3012 & n3020;
  assign n3022 =  a[30]  & n74;
  assign n3023 =  a[31]  & n3022;
  assign n3024 = ~n587 & n3023;
  assign n3025 =  a[30]  & ~ a[31] ;
  assign n3026 = ~ a[30]  &  a[31] ;
  assign n3027 = ~n3025 & ~n3026;
  assign n3028 = n74 & ~n3027;
  assign n3029 = ~n392 & n3028;
  assign n3030 = ~n3024 & ~n3029;
  assign n3031 = ~n3021 & n3030;
  assign n3032 = ~n3019 & n3031;
  assign n3033 = ~n275 & n2760;
  assign n3034 = ~n292 & n3033;
  assign n3035 = ~n357 & n3034;
  assign n3036 = ~n274 & n3035;
  assign n3037 = ~n245 & n3036;
  assign n3038 = ~n623 & n3037;
  assign n3039 = ~n489 & n3038;
  assign n3040 = ~n286 & ~n453;
  assign n3041 = ~n325 & ~n1127;
  assign n3042 = ~n188 & ~n656;
  assign n3043 = ~n190 & ~n527;
  assign n3044 = ~n400 & ~n713;
  assign n3045 = ~n191 & n3044;
  assign n3046 = n3043 & n3045;
  assign n3047 = n3042 & n3046;
  assign n3048 = n3041 & n3047;
  assign n3049 = n3040 & n3048;
  assign n3050 = n1781 & n3049;
  assign n3051 = n285 & n3050;
  assign n3052 = n3039 & n3051;
  assign n3053 = n533 & n3052;
  assign n3054 = n1141 & n3053;
  assign n3055 = ~n509 & n3054;
  assign n3056 = ~n667 & n3055;
  assign n3057 = ~n563 & n3056;
  assign n3058 = ~n641 & ~n752;
  assign n3059 = ~n637 & n3058;
  assign n3060 = ~n276 & n3059;
  assign n3061 = ~n397 & n3060;
  assign n3062 = ~n490 & n3061;
  assign n3063 = ~n200 & n3062;
  assign n3064 = ~n161 & n3063;
  assign n3065 = ~n1010 & n3064;
  assign n3066 = ~n1246 & n2633;
  assign n3067 = ~n135 & n3066;
  assign n3068 = ~n562 & n3067;
  assign n3069 = n373 & n573;
  assign n3070 = n1438 & n3069;
  assign n3071 = n3068 & n3070;
  assign n3072 = n494 & n3071;
  assign n3073 = n931 & n3072;
  assign n3074 = n2317 & n3073;
  assign n3075 = n2651 & n3074;
  assign n3076 = n3065 & n3075;
  assign n3077 = n3057 & n3076;
  assign n3078 = n804 & n3077;
  assign n3079 = ~n427 & n3078;
  assign n3080 = ~n353 & n3079;
  assign n3081 = ~n1102 & n3080;
  assign n3082 = ~n203 & n3081;
  assign n3083 = ~n240 & n3082;
  assign n3084 = ~n203 & ~n791;
  assign n3085 = ~n532 & n3084;
  assign n3086 = n723 & n3085;
  assign n3087 = n615 & n3086;
  assign n3088 = ~n1246 & n3087;
  assign n3089 = ~n135 & n3088;
  assign n3090 = ~n328 & n3089;
  assign n3091 = ~n290 & n3090;
  assign n3092 = ~n961 & n3091;
  assign n3093 = ~n142 & n3092;
  assign n3094 = ~n358 & n3093;
  assign n3095 = n497 & n3059;
  assign n3096 = n3094 & n3095;
  assign n3097 = n2698 & n3096;
  assign n3098 = n2573 & n3097;
  assign n3099 = n1827 & n3098;
  assign n3100 = n1884 & n3099;
  assign n3101 = ~n136 & n3100;
  assign n3102 = ~n177 & n3101;
  assign n3103 = ~n118 & n3102;
  assign n3104 = ~n228 & n3103;
  assign n3105 = ~n287 & n3104;
  assign n3106 = ~n505 & n3105;
  assign n3107 = ~n170 & n3106;
  assign n3108 = ~n666 & n3107;
  assign n3109 = ~n462 & n2191;
  assign n3110 = ~n713 & n3109;
  assign n3111 = ~n281 & n3110;
  assign n3112 = ~n173 & n3111;
  assign n3113 = ~n1203 & n3112;
  assign n3114 = ~n275 & n2347;
  assign n3115 = ~n168 & n968;
  assign n3116 = n1333 & n3115;
  assign n3117 = n3114 & n3116;
  assign n3118 = n1132 & n3117;
  assign n3119 = n3113 & n3118;
  assign n3120 = n1917 & n3119;
  assign n3121 = n2678 & n3120;
  assign n3122 = n1781 & n3121;
  assign n3123 = n1366 & n3122;
  assign n3124 = n1248 & n3123;
  assign n3125 = ~n242 & n3124;
  assign n3126 = ~n191 & n3125;
  assign n3127 = ~n127 & n3126;
  assign n3128 = n618 & ~n847;
  assign n3129 = n897 & n3128;
  assign n3130 = n439 & n3129;
  assign n3131 = n690 & n3130;
  assign n3132 = n2091 & n3131;
  assign n3133 = n1126 & n3132;
  assign n3134 = n1488 & n3133;
  assign n3135 = n3127 & n3134;
  assign n3136 = n512 & n3135;
  assign n3137 = n3108 & n3136;
  assign n3138 = n1994 & n3137;
  assign n3139 = n1237 & n3138;
  assign n3140 = n341 & n3139;
  assign n3141 = ~n1306 & n3140;
  assign n3142 = ~n461 & n3141;
  assign n3143 = ~n403 & n3142;
  assign n3144 = ~n492 & n3143;
  assign n3145 = ~n163 & n3144;
  assign n3146 = ~n271 & n3145;
  assign n3147 = ~n334 & ~n462;
  assign n3148 = ~n531 & n3147;
  assign n3149 = n128 & n3148;
  assign n3150 = n2467 & n3149;
  assign n3151 = ~n505 & n3150;
  assign n3152 = ~n466 & n3151;
  assign n3153 = ~n519 & n3152;
  assign n3154 = ~n251 & n3153;
  assign n3155 = ~n363 & n3154;
  assign n3156 = n876 & n2808;
  assign n3157 = ~n402 & n3156;
  assign n3158 = ~n460 & n3157;
  assign n3159 = ~n298 & n3158;
  assign n3160 = ~n325 & ~n803;
  assign n3161 = ~n712 & n747;
  assign n3162 = ~n1010 & n3161;
  assign n3163 = ~n168 & ~n425;
  assign n3164 = ~n474 & n3163;
  assign n3165 = ~n222 & n3164;
  assign n3166 = n2349 & n3165;
  assign n3167 = n3162 & n3166;
  assign n3168 = n3160 & n3167;
  assign n3169 = n665 & n3168;
  assign n3170 = n2633 & n3169;
  assign n3171 = n1063 & n3170;
  assign n3172 = n1139 & n3171;
  assign n3173 = n804 & n3172;
  assign n3174 = n3159 & n3173;
  assign n3175 = n810 & n3174;
  assign n3176 = n341 & n3175;
  assign n3177 = ~n136 & n3176;
  assign n3178 = ~n255 & n3177;
  assign n3179 = ~n656 & n3178;
  assign n3180 = ~n417 & n3179;
  assign n3181 = n401 & n510;
  assign n3182 = n193 & n3181;
  assign n3183 = ~n111 & n3182;
  assign n3184 = ~n203 & n3183;
  assign n3185 = ~n368 & n3184;
  assign n3186 = ~n163 & n3185;
  assign n3187 = ~n273 & n3186;
  assign n3188 = ~n237 & n3187;
  assign n3189 = ~n225 & n3188;
  assign n3190 = ~n295 & n3189;
  assign n3191 = ~n270 & n3190;
  assign n3192 = n507 & ~n1011;
  assign n3193 = ~n276 & ~n330;
  assign n3194 = ~n152 & n3193;
  assign n3195 = n3192 & n3194;
  assign n3196 = n1423 & n3195;
  assign n3197 = n1555 & n3196;
  assign n3198 = n3191 & n3197;
  assign n3199 = n1825 & n3198;
  assign n3200 = n731 & n3199;
  assign n3201 = n1252 & n3200;
  assign n3202 = ~n514 & n3201;
  assign n3203 = ~n327 & n3202;
  assign n3204 = ~n142 & n3203;
  assign n3205 = ~n99 & n3204;
  assign n3206 = ~n224 & ~n329;
  assign n3207 = ~n617 & n3206;
  assign n3208 = ~n236 & n3207;
  assign n3209 = ~n420 & n3208;
  assign n3210 = ~n752 & n3209;
  assign n3211 = ~n1101 & n3210;
  assign n3212 = ~n248 & n3211;
  assign n3213 = ~n102 & n3212;
  assign n3214 = ~n825 & n3213;
  assign n3215 = ~n167 & n3214;
  assign n3216 = ~n791 & n3215;
  assign n3217 = ~n338 & n3216;
  assign n3218 = ~n592 & n3217;
  assign n3219 = ~n188 & n3218;
  assign n3220 = n674 & n1531;
  assign n3221 = ~n130 & n3220;
  assign n3222 = ~n468 & n3221;
  assign n3223 = ~n1127 & n3222;
  assign n3224 = ~n95 & n3223;
  assign n3225 = ~n429 & n3224;
  assign n3226 = ~n233 & ~n395;
  assign n3227 = n2332 & n3226;
  assign n3228 = n3225 & n3227;
  assign n3229 = n3219 & n3228;
  assign n3230 = n3205 & n3229;
  assign n3231 = n3180 & n3230;
  assign n3232 = n3155 & n3231;
  assign n3233 = n120 & n3232;
  assign n3234 = n621 & n3233;
  assign n3235 = n1574 & n3234;
  assign n3236 = ~n713 & n3235;
  assign n3237 = ~n358 & n3236;
  assign n3238 = ~n158 & n3237;
  assign n3239 = ~n249 & n3238;
  assign n3240 = ~n3146 & ~n3239;
  assign n3241 = n3146 & n3239;
  assign n3242 = ~n3240 & ~n3241;
  assign n3243 = ~ a[20]  & n3242;
  assign n3244 = ~n3240 & ~n3243;
  assign n3245 = n3083 & ~n3244;
  assign n3246 = ~n3083 & n3244;
  assign n3247 = ~n3245 & ~n3246;
  assign n3248 = ~n3032 & n3247;
  assign n3249 = ~n3032 & ~n3248;
  assign n3250 = n3247 & ~n3248;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = ~n173 & ~n226;
  assign n3253 = ~n398 & n2705;
  assign n3254 = ~n154 & n3253;
  assign n3255 = ~n281 & n3254;
  assign n3256 = ~n656 & n3255;
  assign n3257 = ~n637 & n3256;
  assign n3258 = ~n192 & n3257;
  assign n3259 = ~n791 & n3258;
  assign n3260 = ~n255 & n1394;
  assign n3261 = ~n273 & n3260;
  assign n3262 = ~n354 & n539;
  assign n3263 = ~n224 & n3262;
  assign n3264 = ~n666 & n3263;
  assign n3265 = ~n271 & n471;
  assign n3266 = ~n363 & n3265;
  assign n3267 = n1063 & n1128;
  assign n3268 = ~n225 & n3267;
  assign n3269 = n3266 & n3268;
  assign n3270 = n3264 & n3269;
  assign n3271 = n2931 & n3270;
  assign n3272 = n1012 & n3271;
  assign n3273 = n3261 & n3272;
  assign n3274 = n3259 & n3273;
  assign n3275 = n773 & n3274;
  assign n3276 = n291 & n3275;
  assign n3277 = ~n353 & n3276;
  assign n3278 = ~n641 & n3277;
  assign n3279 = ~n352 & n3278;
  assign n3280 = ~n563 & n3279;
  assign n3281 = ~n633 & n3280;
  assign n3282 = ~n188 & n3281;
  assign n3283 = ~n557 & ~n1246;
  assign n3284 = ~n803 & n3283;
  assign n3285 = ~n334 & n3284;
  assign n3286 = ~n299 & n3285;
  assign n3287 = ~n527 & n3286;
  assign n3288 = ~n639 & n3287;
  assign n3289 = ~n525 & n3288;
  assign n3290 = ~n270 & n3289;
  assign n3291 = ~n280 & n720;
  assign n3292 = ~n715 & n3291;
  assign n3293 = ~n961 & n3292;
  assign n3294 = ~n142 & n3293;
  assign n3295 = ~n932 & n3294;
  assign n3296 = ~n531 & n3295;
  assign n3297 = ~n205 & n2651;
  assign n3298 = ~n222 & n3297;
  assign n3299 = ~n395 & ~n452;
  assign n3300 = ~n489 & n3299;
  assign n3301 = n3298 & n3300;
  assign n3302 = n3296 & n3301;
  assign n3303 = n1523 & n3302;
  assign n3304 = n3290 & n3303;
  assign n3305 = n1479 & n3304;
  assign n3306 = n128 & n3305;
  assign n3307 = n423 & n3306;
  assign n3308 = n731 & n3307;
  assign n3309 = n507 & n3308;
  assign n3310 = ~n393 & n3309;
  assign n3311 = ~n451 & n3310;
  assign n3312 = ~n231 & n3311;
  assign n3313 = ~n397 & ~n435;
  assign n3314 = ~n438 & n3313;
  assign n3315 = n1071 & n3314;
  assign n3316 = n1931 & n3315;
  assign n3317 = n524 & n3316;
  assign n3318 = n2237 & n3317;
  assign n3319 = n3312 & n3318;
  assign n3320 = n3282 & n3319;
  assign n3321 = n872 & n3320;
  assign n3322 = n3252 & n3321;
  assign n3323 = n804 & n3322;
  assign n3324 = n570 & n3323;
  assign n3325 = ~n233 & n3324;
  assign n3326 = ~n594 & n3325;
  assign n3327 = ~n158 & n3326;
  assign n3328 = n3146 & ~n3327;
  assign n3329 = ~n3146 & n3327;
  assign n3330 = n2920 & ~n2922;
  assign n3331 = ~n2923 & ~n3330;
  assign n3332 = n75 & n3331;
  assign n3333 = ~n587 & n3020;
  assign n3334 = ~n867 & n3023;
  assign n3335 = ~n710 & n3028;
  assign n3336 = ~n3334 & ~n3335;
  assign n3337 = ~n3333 & n3336;
  assign n3338 = ~n3332 & n3337;
  assign n3339 = ~n3328 & ~n3338;
  assign n3340 = ~n3329 & n3339;
  assign n3341 = ~n3328 & ~n3340;
  assign n3342 = ~ a[20]  & ~n3243;
  assign n3343 = ~n3241 & n3244;
  assign n3344 = ~n3342 & ~n3343;
  assign n3345 = ~n3341 & ~n3344;
  assign n3346 = n2924 & ~n2926;
  assign n3347 = ~n2927 & ~n3346;
  assign n3348 = n75 & n3347;
  assign n3349 = ~n392 & n3020;
  assign n3350 = ~n710 & n3023;
  assign n3351 = ~n587 & n3028;
  assign n3352 = ~n3350 & ~n3351;
  assign n3353 = ~n3349 & n3352;
  assign n3354 = ~n3348 & n3353;
  assign n3355 = n3341 & n3344;
  assign n3356 = ~n3345 & ~n3355;
  assign n3357 = ~n3354 & n3356;
  assign n3358 = ~n3345 & ~n3357;
  assign n3359 = ~n3251 & ~n3358;
  assign n3360 = n3251 & n3358;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 =  a[28]  & ~ a[29] ;
  assign n3363 = ~ a[28]  &  a[29] ;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 =  a[26]  & ~ a[27] ;
  assign n3366 = ~ a[26]  &  a[27] ;
  assign n3367 = ~n3365 & ~n3366;
  assign n3368 = ~n3364 & ~n3367;
  assign n3369 = ~n469 & ~n656;
  assign n3370 = ~n1010 & n3369;
  assign n3371 = n2426 & n3370;
  assign n3372 = n2361 & n3371;
  assign n3373 = ~n194 & n3372;
  assign n3374 = ~n746 & n3373;
  assign n3375 = ~n339 & n3374;
  assign n3376 = ~n145 & n3375;
  assign n3377 = ~n567 & n3376;
  assign n3378 = ~n393 & n3377;
  assign n3379 = ~n146 & ~n536;
  assign n3380 = ~n428 & n3379;
  assign n3381 = ~n301 & n3380;
  assign n3382 = ~n511 & n3381;
  assign n3383 = ~n461 & n3382;
  assign n3384 = ~n563 & n3383;
  assign n3385 = ~n689 & n3384;
  assign n3386 = ~n200 & n3385;
  assign n3387 = ~n1306 & n2508;
  assign n3388 = ~n154 & n3387;
  assign n3389 = ~n417 & n3388;
  assign n3390 = ~n372 & ~n427;
  assign n3391 = ~n332 & n3390;
  assign n3392 = n937 & n1181;
  assign n3393 = ~n641 & n3392;
  assign n3394 = n1392 & n1739;
  assign n3395 = n3393 & n3394;
  assign n3396 = n3391 & n3395;
  assign n3397 = n3389 & n3396;
  assign n3398 = n3386 & n3397;
  assign n3399 = n291 & n3398;
  assign n3400 = ~n617 & n3399;
  assign n3401 = ~n135 & n3400;
  assign n3402 = ~n460 & n3401;
  assign n3403 = ~n451 & n3402;
  assign n3404 = ~n337 & n3403;
  assign n3405 = ~n875 & n3404;
  assign n3406 = ~n667 & n2073;
  assign n3407 = ~n752 & n3406;
  assign n3408 = ~n118 & n3407;
  assign n3409 = ~n254 & ~n335;
  assign n3410 = n300 & n962;
  assign n3411 = n3409 & n3410;
  assign n3412 = ~n1072 & n3411;
  assign n3413 = ~n513 & n3412;
  assign n3414 = ~n191 & n3413;
  assign n3415 = ~n712 & n3414;
  assign n3416 = n116 & n515;
  assign n3417 = n1045 & n3416;
  assign n3418 = n3266 & n3417;
  assign n3419 = n1388 & n3418;
  assign n3420 = n1132 & n3419;
  assign n3421 = n3415 & n3420;
  assign n3422 = n3408 & n3421;
  assign n3423 = n1528 & n3422;
  assign n3424 = n873 & n3423;
  assign n3425 = n1182 & n3424;
  assign n3426 = n720 & n3425;
  assign n3427 = ~n121 & n3426;
  assign n3428 = ~n305 & n3427;
  assign n3429 = ~n226 & n3428;
  assign n3430 = ~n403 & n3429;
  assign n3431 = ~n206 & n3430;
  assign n3432 = ~n492 & n3431;
  assign n3433 = ~n352 & n1141;
  assign n3434 = ~n537 & n3433;
  assign n3435 = ~n603 & n3434;
  assign n3436 = ~n568 & ~n716;
  assign n3437 = ~n142 & n3436;
  assign n3438 = ~n86 & ~n240;
  assign n3439 = n3437 & n3438;
  assign n3440 = n3435 & n3439;
  assign n3441 = n3225 & n3440;
  assign n3442 = n3432 & n3441;
  assign n3443 = n3405 & n3442;
  assign n3444 = n2740 & n3443;
  assign n3445 = n3378 & n3444;
  assign n3446 = n247 & n3445;
  assign n3447 = n1917 & n3446;
  assign n3448 = n491 & n3447;
  assign n3449 = n978 & n3448;
  assign n3450 = n810 & n3449;
  assign n3451 = ~n462 & n3450;
  assign n3452 = ~n777 & n3451;
  assign n3453 = ~n225 & n3452;
  assign n3454 = ~n304 & n3453;
  assign n3455 = ~n295 & n3454;
  assign n3456 = ~n519 & n3455;
  assign n3457 = n3364 & ~n3367;
  assign n3458 = ~n3456 & n3457;
  assign n3459 = ~n119 & ~n271;
  assign n3460 = ~n254 & n3459;
  assign n3461 = ~n496 & n3460;
  assign n3462 = ~n536 & n3461;
  assign n3463 = ~n712 & n3462;
  assign n3464 = ~n1010 & n3463;
  assign n3465 = n792 & n2091;
  assign n3466 = ~n1101 & n3465;
  assign n3467 = ~n296 & n3466;
  assign n3468 = ~n980 & n3467;
  assign n3469 = ~n623 & n3468;
  assign n3470 = ~n525 & n3469;
  assign n3471 = ~n331 & n2105;
  assign n3472 = ~n453 & n3471;
  assign n3473 = n418 & ~n469;
  assign n3474 = ~n474 & n3473;
  assign n3475 = n754 & n3226;
  assign n3476 = n3474 & n3475;
  assign n3477 = n2556 & n3476;
  assign n3478 = n593 & n3477;
  assign n3479 = n437 & n3478;
  assign n3480 = n1601 & n3479;
  assign n3481 = n3472 & n3480;
  assign n3482 = n615 & n3481;
  assign n3483 = n1046 & n3482;
  assign n3484 = n3470 & n3483;
  assign n3485 = n1576 & n3484;
  assign n3486 = n570 & n3485;
  assign n3487 = ~n330 & n3486;
  assign n3488 = ~n302 & n3487;
  assign n3489 = ~n164 & n3488;
  assign n3490 = ~n157 & ~n571;
  assign n3491 = n401 & n2113;
  assign n3492 = n1531 & n3491;
  assign n3493 = ~n355 & n3492;
  assign n3494 = ~n284 & n3493;
  assign n3495 = ~n777 & n3494;
  assign n3496 = ~n206 & n3495;
  assign n3497 = ~n237 & n3496;
  assign n3498 = n941 & n1255;
  assign n3499 = n2220 & n3498;
  assign n3500 = n2007 & n3499;
  assign n3501 = n3497 & n3500;
  assign n3502 = n614 & n3501;
  assign n3503 = n2021 & n3502;
  assign n3504 = n291 & n3503;
  assign n3505 = n1269 & n3504;
  assign n3506 = ~n617 & n3505;
  assign n3507 = ~n224 & n3506;
  assign n3508 = ~n419 & n3507;
  assign n3509 = n3490 & n3508;
  assign n3510 = ~n366 & n3509;
  assign n3511 = ~n248 & ~n426;
  assign n3512 = ~n715 & n3511;
  assign n3513 = n968 & ~n1062;
  assign n3514 = ~n425 & n3513;
  assign n3515 = n172 & n3514;
  assign n3516 = n3512 & n3515;
  assign n3517 = n2022 & n3516;
  assign n3518 = n3510 & n3517;
  assign n3519 = ~n847 & n3518;
  assign n3520 = ~n961 & n3519;
  assign n3521 = ~n245 & n3520;
  assign n3522 = ~n121 & ~n145;
  assign n3523 = ~n338 & n3522;
  assign n3524 = ~n286 & ~n332;
  assign n3525 = n3298 & n3524;
  assign n3526 = n3523 & n3525;
  assign n3527 = n530 & n3526;
  assign n3528 = n1586 & n3527;
  assign n3529 = n465 & n3528;
  assign n3530 = n3521 & n3529;
  assign n3531 = n3489 & n3530;
  assign n3532 = n3464 & n3531;
  assign n3533 = n1029 & n3532;
  assign n3534 = n1528 & n3533;
  assign n3535 = n1254 & n3534;
  assign n3536 = n591 & n3535;
  assign n3537 = ~n334 & n3536;
  assign n3538 = ~n192 & n3537;
  assign n3539 = ~n371 & n3538;
  assign n3540 = ~n79 & ~n82;
  assign n3541 = ~n3364 & n3367;
  assign n3542 = ~n3540 & n3541;
  assign n3543 = ~n3539 & n3542;
  assign n3544 = ~n233 & ~n884;
  assign n3545 = ~n713 & ~n791;
  assign n3546 = ~n375 & n3545;
  assign n3547 = ~n332 & n3546;
  assign n3548 = ~n569 & n3547;
  assign n3549 = ~n226 & ~n1127;
  assign n3550 = n1960 & n3549;
  assign n3551 = n3548 & n3550;
  assign n3552 = n2010 & n3551;
  assign n3553 = n1479 & n3552;
  assign n3554 = n3544 & n3553;
  assign n3555 = n1574 & n3554;
  assign n3556 = n421 & n3555;
  assign n3557 = ~n354 & n3556;
  assign n3558 = ~n334 & n3557;
  assign n3559 = ~n623 & n3558;
  assign n3560 = n116 & ~n1306;
  assign n3561 = ~n506 & n3560;
  assign n3562 = ~n326 & n3561;
  assign n3563 = ~n568 & n3562;
  assign n3564 = ~n430 & n3563;
  assign n3565 = ~n422 & n3564;
  assign n3566 = ~n495 & ~n619;
  assign n3567 = ~n357 & n3566;
  assign n3568 = ~n777 & n3567;
  assign n3569 = ~n490 & n3568;
  assign n3570 = ~n428 & n2582;
  assign n3571 = n2267 & n3570;
  assign n3572 = n2013 & n3571;
  assign n3573 = n2348 & n3572;
  assign n3574 = n3569 & n3573;
  assign n3575 = ~n462 & n3574;
  assign n3576 = ~n563 & n3575;
  assign n3577 = ~n536 & n3576;
  assign n3578 = ~n132 & n3577;
  assign n3579 = ~n338 & n3578;
  assign n3580 = ~n337 & n3579;
  assign n3581 = ~n355 & ~n426;
  assign n3582 = ~n396 & n3581;
  assign n3583 = ~n470 & n3582;
  assign n3584 = n1330 & n1826;
  assign n3585 = ~n398 & n3584;
  assign n3586 = ~n95 & n3585;
  assign n3587 = ~n358 & n3586;
  assign n3588 = n3583 & n3587;
  assign n3589 = n3580 & n3588;
  assign n3590 = n1928 & n3589;
  assign n3591 = n3565 & n3590;
  assign n3592 = n221 & n3591;
  assign n3593 = n1687 & n3592;
  assign n3594 = n3559 & n3593;
  assign n3595 = ~n236 & n3594;
  assign n3596 = ~n135 & n3595;
  assign n3597 = ~n280 & n3596;
  assign n3598 = ~n1101 & n3597;
  assign n3599 = ~n514 & n3598;
  assign n3600 = ~n305 & n3599;
  assign n3601 = ~n689 & n3600;
  assign n3602 = ~n304 & n3601;
  assign n3603 = ~n86 & n3602;
  assign n3604 = ~n489 & n3603;
  assign n3605 = ~n771 & n3604;
  assign n3606 = n3367 & n3540;
  assign n3607 = ~n3605 & n3606;
  assign n3608 = ~n3543 & ~n3607;
  assign n3609 = ~n3458 & n3608;
  assign n3610 = ~n3368 & n3609;
  assign n3611 = ~n3539 & ~n3605;
  assign n3612 = ~n3012 & ~n3539;
  assign n3613 = ~n3013 & ~n3016;
  assign n3614 = n3012 & n3539;
  assign n3615 = ~n3612 & ~n3614;
  assign n3616 = ~n3613 & n3615;
  assign n3617 = ~n3612 & ~n3616;
  assign n3618 = n3539 & n3605;
  assign n3619 = ~n3611 & ~n3618;
  assign n3620 = ~n3617 & n3619;
  assign n3621 = ~n3611 & ~n3620;
  assign n3622 = ~n3456 & ~n3605;
  assign n3623 = n3456 & n3605;
  assign n3624 = ~n3622 & ~n3623;
  assign n3625 = ~n3621 & n3624;
  assign n3626 = n3621 & ~n3624;
  assign n3627 = ~n3625 & ~n3626;
  assign n3628 = n3609 & ~n3627;
  assign n3629 = ~n3610 & ~n3628;
  assign n3630 =  a[29]  & ~n3629;
  assign n3631 = ~ a[29]  & n3629;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = n3361 & ~n3632;
  assign n3634 = ~n3359 & ~n3633;
  assign n3635 = ~n3245 & ~n3248;
  assign n3636 = ~n619 & n1531;
  assign n3637 = ~n509 & n3226;
  assign n3638 = ~n511 & n3637;
  assign n3639 = ~n1062 & n3638;
  assign n3640 = ~n656 & n3639;
  assign n3641 = ~n149 & n3640;
  assign n3642 = ~n367 & n3641;
  assign n3643 = ~n245 & n3642;
  assign n3644 = ~n81 & n3643;
  assign n3645 = ~n132 & ~n163;
  assign n3646 = n202 & n3645;
  assign n3647 = ~n557 & n3646;
  assign n3648 = ~n353 & n3647;
  assign n3649 = ~n175 & n3648;
  assign n3650 = ~n243 & n3649;
  assign n3651 = ~n569 & n3650;
  assign n3652 = n1408 & n1458;
  assign n3653 = n3472 & n3652;
  assign n3654 = n3252 & n3653;
  assign n3655 = ~n398 & n3654;
  assign n3656 = ~n232 & n3655;
  assign n3657 = ~n171 & n3656;
  assign n3658 = ~n299 & n3657;
  assign n3659 = ~n357 & n3658;
  assign n3660 = ~n374 & n3659;
  assign n3661 = ~n368 & n3660;
  assign n3662 = ~n95 & n3661;
  assign n3663 = ~n633 & n3662;
  assign n3664 = n3651 & n3663;
  assign n3665 = n2581 & n3664;
  assign n3666 = n3644 & n3665;
  assign n3667 = n241 & n3666;
  assign n3668 = ~n136 & n3667;
  assign n3669 = n3636 & n3668;
  assign n3670 = ~n425 & n3669;
  assign n3671 = ~n274 & n3670;
  assign n3672 = ~n466 & n3671;
  assign n3673 = ~n422 & n3672;
  assign n3674 = ~n338 & n3673;
  assign n3675 = ~n655 & n3674;
  assign n3676 = ~n229 & ~n1072;
  assign n3677 = ~n275 & n3676;
  assign n3678 = ~n461 & n3677;
  assign n3679 = ~n416 & n3678;
  assign n3680 = ~n1203 & n3679;
  assign n3681 = ~n252 & n3680;
  assign n3682 = ~n504 & ~n641;
  assign n3683 = ~n306 & n3682;
  assign n3684 = ~n272 & n3683;
  assign n3685 = ~n222 & n3684;
  assign n3686 = ~n493 & n1380;
  assign n3687 = ~n1010 & n3686;
  assign n3688 = n2427 & n3687;
  assign n3689 = n723 & n3688;
  assign n3690 = n3685 & n3689;
  assign n3691 = n1323 & n3690;
  assign n3692 = n3681 & n3691;
  assign n3693 = n3675 & n3692;
  assign n3694 = n1915 & n3693;
  assign n3695 = n1046 & n3694;
  assign n3696 = n1366 & n3695;
  assign n3697 = ~n169 & n3696;
  assign n3698 = ~n847 & n3697;
  assign n3699 = ~n151 & n3698;
  assign n3700 = ~n118 & n3699;
  assign n3701 = ~n206 & n3700;
  assign n3702 = ~n452 & n3701;
  assign n3703 = n3083 & ~n3702;
  assign n3704 = ~n3083 & n3702;
  assign n3705 = ~n3635 & ~n3704;
  assign n3706 = ~n3703 & n3705;
  assign n3707 = ~n3635 & ~n3706;
  assign n3708 = ~n3704 & ~n3706;
  assign n3709 = ~n3703 & n3708;
  assign n3710 = ~n3707 & ~n3709;
  assign n3711 = n3020 & ~n3539;
  assign n3712 = ~n3012 & n3028;
  assign n3713 = ~n392 & n3023;
  assign n3714 = n3613 & ~n3615;
  assign n3715 = ~n3616 & ~n3714;
  assign n3716 = n75 & n3715;
  assign n3717 = ~n3713 & ~n3716;
  assign n3718 = ~n3712 & n3717;
  assign n3719 = ~n3711 & n3718;
  assign n3720 = ~n3710 & ~n3719;
  assign n3721 = ~n3710 & ~n3720;
  assign n3722 = ~n3719 & ~n3720;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3634 & ~n3723;
  assign n3725 = ~n3634 & ~n3724;
  assign n3726 = ~n3723 & ~n3724;
  assign n3727 = ~n3725 & ~n3726;
  assign n3728 = ~n189 & ~n280;
  assign n3729 = ~n115 & n3728;
  assign n3730 = ~n169 & n3729;
  assign n3731 = ~n149 & n3730;
  assign n3732 = ~n490 & n3731;
  assign n3733 = ~n567 & n3732;
  assign n3734 = ~n558 & n1839;
  assign n3735 = ~n667 & n3734;
  assign n3736 = ~n752 & n3735;
  assign n3737 = ~n557 & n3736;
  assign n3738 = ~n223 & n3737;
  assign n3739 = ~n623 & n3738;
  assign n3740 = n640 & n895;
  assign n3741 = ~n123 & n3740;
  assign n3742 = ~n150 & n3741;
  assign n3743 = ~n231 & n3742;
  assign n3744 = n401 & n2556;
  assign n3745 = n3743 & n3744;
  assign n3746 = n3739 & n3745;
  assign n3747 = n3733 & n3746;
  assign n3748 = n2582 & n3747;
  assign n3749 = n720 & n3748;
  assign n3750 = n1141 & n3749;
  assign n3751 = n515 & n3750;
  assign n3752 = n1367 & n3751;
  assign n3753 = ~n803 & n3752;
  assign n3754 = ~n511 & n3753;
  assign n3755 = ~n177 & n3754;
  assign n3756 = ~n147 & n3755;
  assign n3757 = ~n425 & n3756;
  assign n3758 = ~n620 & n2293;
  assign n3759 = ~n205 & n3758;
  assign n3760 = ~n161 & n3759;
  assign n3761 = ~n474 & n3760;
  assign n3762 = ~n340 & n3761;
  assign n3763 = ~n436 & n3762;
  assign n3764 = ~n564 & n3763;
  assign n3765 = n1392 & n3115;
  assign n3766 = n590 & n3765;
  assign n3767 = ~n118 & n3766;
  assign n3768 = ~n527 & n3767;
  assign n3769 = ~n422 & n747;
  assign n3770 = ~n1010 & n3769;
  assign n3771 = ~n569 & n3770;
  assign n3772 = n1784 & n3771;
  assign n3773 = n3768 & n3772;
  assign n3774 = n2512 & n3773;
  assign n3775 = n872 & n3774;
  assign n3776 = ~n276 & n3775;
  assign n3777 = ~n602 & n3776;
  assign n3778 = ~n884 & n3777;
  assign n3779 = ~n394 & n3778;
  assign n3780 = ~n325 & n3779;
  assign n3781 = ~n271 & n3780;
  assign n3782 = ~n428 & n3781;
  assign n3783 = n1388 & n1577;
  assign n3784 = ~n563 & n3783;
  assign n3785 = ~n132 & n3784;
  assign n3786 = ~n225 & n3785;
  assign n3787 = ~n531 & n3786;
  assign n3788 = ~n657 & n3787;
  assign n3789 = ~n1104 & n3788;
  assign n3790 = ~n86 & n3789;
  assign n3791 = ~n144 & ~n466;
  assign n3792 = ~n191 & n3791;
  assign n3793 = n3040 & n3792;
  assign n3794 = n3790 & n3793;
  assign n3795 = n3782 & n3794;
  assign n3796 = n3764 & n3795;
  assign n3797 = n2740 & n3796;
  assign n3798 = n937 & n3797;
  assign n3799 = n3757 & n3798;
  assign n3800 = n1761 & n3799;
  assign n3801 = n538 & n3800;
  assign n3802 = ~n462 & n3801;
  assign n3803 = ~n402 & n3802;
  assign n3804 = ~n277 & n3803;
  assign n3805 = ~n293 & n3804;
  assign n3806 = n3457 & ~n3805;
  assign n3807 = n3542 & ~n3605;
  assign n3808 = ~n3456 & n3606;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = ~n3806 & n3809;
  assign n3811 = ~n3368 & n3810;
  assign n3812 = ~n3622 & ~n3625;
  assign n3813 = ~n3456 & ~n3805;
  assign n3814 = n3456 & n3805;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = ~n3812 & n3815;
  assign n3817 = n3812 & ~n3815;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = n3810 & ~n3818;
  assign n3820 = ~n3811 & ~n3819;
  assign n3821 =  a[29]  & ~n3820;
  assign n3822 = ~ a[29]  & n3820;
  assign n3823 = ~n3821 & ~n3822;
  assign n3824 = n3727 & n3823;
  assign n3825 = ~n3727 & ~n3823;
  assign n3826 = ~n3824 & ~n3825;
  assign n3827 = ~n286 & ~n438;
  assign n3828 = n3437 & n3827;
  assign n3829 = ~n245 & n3828;
  assign n3830 = ~n791 & n3829;
  assign n3831 = ~n422 & n3830;
  assign n3832 = ~n298 & ~n961;
  assign n3833 = n3831 & n3832;
  assign n3834 = n665 & n3833;
  assign n3835 = n539 & n3834;
  assign n3836 = n454 & n3835;
  assign n3837 = n193 & n3836;
  assign n3838 = ~n99 & n3837;
  assign n3839 = ~n372 & n3838;
  assign n3840 = n772 & n1105;
  assign n3841 = n471 & n3840;
  assign n3842 = n827 & n3841;
  assign n3843 = ~n657 & n3842;
  assign n3844 = ~n252 & n3843;
  assign n3845 = ~n592 & n3844;
  assign n3846 = ~n277 & n3845;
  assign n3847 = ~n332 & n3846;
  assign n3848 = ~n1127 & n3847;
  assign n3849 = n2208 & n2573;
  assign n3850 = n128 & n3849;
  assign n3851 = ~n489 & n3850;
  assign n3852 = ~n119 & n3851;
  assign n3853 = n2275 & n3852;
  assign n3854 = n3848 & n3853;
  assign n3855 = ~n86 & n3854;
  assign n3856 = ~n569 & n3855;
  assign n3857 = ~n429 & n590;
  assign n3858 = ~n231 & n3857;
  assign n3859 = n624 & n3206;
  assign n3860 = n2963 & n3859;
  assign n3861 = n1254 & n3860;
  assign n3862 = n979 & n3861;
  assign n3863 = n356 & n3862;
  assign n3864 = ~n289 & n3863;
  assign n3865 = ~n284 & n3864;
  assign n3866 = ~n557 & n3865;
  assign n3867 = n3858 & n3866;
  assign n3868 = ~n633 & n3867;
  assign n3869 = ~n270 & n3868;
  assign n3870 = n3570 & n3869;
  assign n3871 = n1480 & n3870;
  assign n3872 = n968 & n3871;
  assign n3873 = ~n449 & n3872;
  assign n3874 = n3856 & n3873;
  assign n3875 = n3839 & n3874;
  assign n3876 = ~n328 & n3875;
  assign n3877 = ~n296 & n3876;
  assign n3878 =  a[23]  & ~ a[24] ;
  assign n3879 = ~ a[23]  &  a[24] ;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 =  a[25]  & ~ a[26] ;
  assign n3882 = ~ a[25]  &  a[26] ;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = ~n3880 & n3883;
  assign n3885 = ~n3877 & n3884;
  assign n3886 = ~n127 & ~n277;
  assign n3887 = n2390 & n3041;
  assign n3888 = n2633 & n3887;
  assign n3889 = n1479 & n3888;
  assign n3890 = n1824 & n3889;
  assign n3891 = n3886 & n3890;
  assign n3892 = ~n190 & n3891;
  assign n3893 = ~n847 & n3892;
  assign n3894 = ~n777 & n3893;
  assign n3895 = ~n492 & n3894;
  assign n3896 = ~n163 & n3895;
  assign n3897 = ~n170 & n3896;
  assign n3898 = ~n340 & n3897;
  assign n3899 = ~n672 & n3898;
  assign n3900 = ~n436 & n3899;
  assign n3901 = ~n358 & n3900;
  assign n3902 = ~n111 & ~n505;
  assign n3903 = ~n394 & n3902;
  assign n3904 = ~n375 & n3903;
  assign n3905 = ~n883 & n3904;
  assign n3906 = n747 & n978;
  assign n3907 = ~n236 & ~n301;
  assign n3908 = ~n136 & n3907;
  assign n3909 = ~n469 & n3908;
  assign n3910 = ~n1306 & n3909;
  assign n3911 = ~n397 & n3910;
  assign n3912 = ~n398 & n3911;
  assign n3913 = n775 & n3912;
  assign n3914 = ~n1072 & n3913;
  assign n3915 = n517 & n3914;
  assign n3916 = n3906 & n3915;
  assign n3917 = n732 & n3916;
  assign n3918 = n3905 & n3917;
  assign n3919 = n3901 & n3918;
  assign n3920 = n1731 & n3919;
  assign n3921 = ~n617 & n3920;
  assign n3922 = ~n490 & n3921;
  assign n3923 = ~n425 & n3922;
  assign n3924 = ~n468 & n3923;
  assign n3925 = ~n273 & n3924;
  assign n3926 = ~n295 & n3925;
  assign n3927 = ~n532 & n3926;
  assign n3928 = ~n886 & n3927;
  assign n3929 = ~n569 & n3928;
  assign n3930 = ~n330 & n2738;
  assign n3931 = ~n242 & n3930;
  assign n3932 = n2698 & n3931;
  assign n3933 = ~n504 & n3932;
  assign n3934 = ~n245 & n3933;
  assign n3935 = ~n142 & n3934;
  assign n3936 = ~n791 & n3935;
  assign n3937 = ~n567 & n3936;
  assign n3938 = ~n271 & n3937;
  assign n3939 = ~n771 & n3938;
  assign n3940 = n1440 & n3729;
  assign n3941 = n3409 & n3940;
  assign n3942 = n1292 & n3941;
  assign n3943 = ~n276 & n3942;
  assign n3944 = ~n168 & n3943;
  assign n3945 = ~n426 & n3944;
  assign n3946 = ~n1102 & n3945;
  assign n3947 = ~n511 & n3946;
  assign n3948 = ~n372 & n1480;
  assign n3949 = ~n449 & n3948;
  assign n3950 = n1155 & n3949;
  assign n3951 = n3947 & n3950;
  assign n3952 = n2740 & n3951;
  assign n3953 = n3939 & n3952;
  assign n3954 = n3929 & n3953;
  assign n3955 = n1046 & n3954;
  assign n3956 = n520 & n3955;
  assign n3957 = n2583 & n3956;
  assign n3958 = n720 & n3957;
  assign n3959 = ~n1011 & n3958;
  assign n3960 = ~n980 & n3959;
  assign n3961 = ~n452 & n3960;
  assign n3962 = ~n536 & n3961;
  assign n3963 = ~n283 & n3962;
  assign n3964 = ~n338 & n3963;
  assign n3965 = ~n76 & ~n84;
  assign n3966 = n3880 & ~n3883;
  assign n3967 = ~n3965 & n3966;
  assign n3968 = ~n3964 & n3967;
  assign n3969 = ~n492 & ~n496;
  assign n3970 = ~n430 & n3969;
  assign n3971 = ~n505 & n3970;
  assign n3972 = ~n425 & n3971;
  assign n3973 = n2470 & n3832;
  assign n3974 = ~n619 & n3973;
  assign n3975 = ~n237 & n3974;
  assign n3976 = ~n712 & n3975;
  assign n3977 = ~n451 & n3976;
  assign n3978 = ~n592 & n3977;
  assign n3979 = n1478 & n1726;
  assign n3980 = ~n327 & n3979;
  assign n3981 = ~n91 & n3980;
  assign n3982 = ~n715 & n3981;
  assign n3983 = ~n102 & n3982;
  assign n3984 = ~n287 & n3983;
  assign n3985 = ~n290 & ~n884;
  assign n3986 = ~n147 & n3985;
  assign n3987 = ~n403 & n3986;
  assign n3988 = n1347 & n3987;
  assign n3989 = ~n155 & n3988;
  assign n3990 = ~n396 & n3989;
  assign n3991 = n1916 & n2297;
  assign n3992 = ~n149 & n3991;
  assign n3993 = ~n594 & n3992;
  assign n3994 = ~n223 & n3993;
  assign n3995 = ~n402 & n3994;
  assign n3996 = ~n305 & n3995;
  assign n3997 = ~n226 & n3996;
  assign n3998 = n3990 & n3997;
  assign n3999 = n538 & n3998;
  assign n4000 = ~n435 & n3999;
  assign n4001 = ~n292 & n4000;
  assign n4002 = ~n283 & n4001;
  assign n4003 = ~n372 & n4002;
  assign n4004 = n2133 & n2703;
  assign n4005 = n2739 & n4004;
  assign n4006 = n1248 & n4005;
  assign n4007 = n1389 & n4006;
  assign n4008 = ~n506 & n4007;
  assign n4009 = ~n107 & n4008;
  assign n4010 = ~n275 & n2993;
  assign n4011 = ~n417 & n4010;
  assign n4012 = n3408 & n4011;
  assign n4013 = n4009 & n4012;
  assign n4014 = n4003 & n4013;
  assign n4015 = n1783 & n4014;
  assign n4016 = n421 & n4015;
  assign n4017 = ~n453 & n4016;
  assign n4018 = n3914 & n3931;
  assign n4019 = n3128 & n4018;
  assign n4020 = n3947 & n4019;
  assign n4021 = ~n123 & n4020;
  assign n4022 = ~n194 & n4021;
  assign n4023 = ~n111 & n4022;
  assign n4024 = ~n746 & n4023;
  assign n4025 = ~n462 & n4024;
  assign n4026 = ~n509 & n4025;
  assign n4027 = ~n1011 & n4026;
  assign n4028 = ~n190 & n4027;
  assign n4029 = ~n518 & n4028;
  assign n4030 = ~n151 & n4029;
  assign n4031 = n4017 & n4030;
  assign n4032 = n3984 & n4031;
  assign n4033 = ~n825 & n4032;
  assign n4034 = ~n99 & n4033;
  assign n4035 = n1204 & n3852;
  assign n4036 = n3790 & n4035;
  assign n4037 = n604 & n4036;
  assign n4038 = n1046 & n4037;
  assign n4039 = n159 & n4038;
  assign n4040 = ~n130 & n4039;
  assign n4041 = n4034 & n4040;
  assign n4042 = n3978 & n4041;
  assign n4043 = n3972 & n4042;
  assign n4044 = n471 & n4043;
  assign n4045 = ~n589 & n4044;
  assign n4046 = n3880 & n3965;
  assign n4047 = ~n4045 & n4046;
  assign n4048 = ~n3968 & ~n4047;
  assign n4049 = ~n3885 & n4048;
  assign n4050 = ~n3880 & ~n3883;
  assign n4051 = ~n3964 & ~n4045;
  assign n4052 = ~n3805 & ~n3964;
  assign n4053 = ~n3813 & ~n3816;
  assign n4054 = n3805 & n3964;
  assign n4055 = ~n4052 & ~n4054;
  assign n4056 = ~n4053 & n4055;
  assign n4057 = ~n4052 & ~n4056;
  assign n4058 = n3964 & n4045;
  assign n4059 = ~n4051 & ~n4058;
  assign n4060 = ~n4057 & n4059;
  assign n4061 = ~n4051 & ~n4060;
  assign n4062 = ~n3877 & ~n4045;
  assign n4063 = n3877 & n4045;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = ~n4061 & n4064;
  assign n4066 = n4061 & ~n4064;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = n4050 & n4067;
  assign n4069 = n4049 & ~n4068;
  assign n4070 =  a[26]  & ~n4069;
  assign n4071 =  a[26]  & ~n4070;
  assign n4072 = ~n4069 & ~n4070;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = n3826 & ~n4073;
  assign n4075 = n3826 & ~n4074;
  assign n4076 = ~n4073 & ~n4074;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = n3457 & ~n3605;
  assign n4079 = ~n3012 & n3542;
  assign n4080 = ~n3539 & n3606;
  assign n4081 = ~n4079 & ~n4080;
  assign n4082 = ~n4078 & n4081;
  assign n4083 = n3617 & ~n3619;
  assign n4084 = ~n3620 & ~n4083;
  assign n4085 = n3368 & n4084;
  assign n4086 = n4082 & ~n4085;
  assign n4087 =  a[29]  & ~n4086;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 =  a[29]  & ~n4087;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = ~n3354 & ~n3357;
  assign n4092 = n3356 & ~n3357;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = ~n4090 & ~n4093;
  assign n4095 = ~n4090 & ~n4094;
  assign n4096 = ~n4093 & ~n4094;
  assign n4097 = ~n4095 & ~n4096;
  assign n4098 = ~n3338 & ~n3340;
  assign n4099 = ~n3329 & n3341;
  assign n4100 = ~n4098 & ~n4099;
  assign n4101 = ~n395 & ~n594;
  assign n4102 = ~n354 & ~n1011;
  assign n4103 = ~n177 & n4102;
  assign n4104 = ~n367 & n4103;
  assign n4105 = n250 & n1760;
  assign n4106 = n792 & n4105;
  assign n4107 = n2192 & n4106;
  assign n4108 = n4104 & n4107;
  assign n4109 = n2943 & n4108;
  assign n4110 = n877 & n4109;
  assign n4111 = n2217 & n4110;
  assign n4112 = n3405 & n4111;
  assign n4113 = n3901 & n4112;
  assign n4114 = n2500 & n4113;
  assign n4115 = n1183 & n4114;
  assign n4116 = n507 & n4115;
  assign n4117 = n4101 & n4116;
  assign n4118 = ~n327 & n4117;
  assign n4119 = ~n292 & n4118;
  assign n4120 = ~n286 & n4119;
  assign n4121 = ~n1104 & n4120;
  assign n4122 = ~n395 & n1073;
  assign n4123 = ~n980 & n4122;
  assign n4124 = ~n165 & n4123;
  assign n4125 = ~n932 & n4124;
  assign n4126 = ~n375 & n4125;
  assign n4127 = ~n86 & n4126;
  assign n4128 = n1139 & n1781;
  assign n4129 = ~n242 & n4128;
  assign n4130 = ~n562 & n4129;
  assign n4131 = ~n402 & n1181;
  assign n4132 = ~n416 & n4131;
  assign n4133 = n1045 & n4132;
  assign n4134 = n812 & n4133;
  assign n4135 = n1692 & n4134;
  assign n4136 = n4130 & n4135;
  assign n4137 = n4127 & n4136;
  assign n4138 = n491 & n4137;
  assign n4139 = n1251 & n4138;
  assign n4140 = n1141 & n4139;
  assign n4141 = ~n123 & n4140;
  assign n4142 = ~n334 & n4141;
  assign n4143 = ~n1101 & n4142;
  assign n4144 = ~n594 & n4143;
  assign n4145 = ~n527 & n4144;
  assign n4146 = ~n689 & n4145;
  assign n4147 = ~n200 & n4146;
  assign n4148 = ~n1104 & n4147;
  assign n4149 = ~n168 & ~n1203;
  assign n4150 = ~n886 & n4149;
  assign n4151 = ~n188 & n4150;
  assign n4152 = n279 & ~n589;
  assign n4153 = ~n394 & n4152;
  assign n4154 = n4151 & n4153;
  assign n4155 = n2371 & n4154;
  assign n4156 = n3521 & n4155;
  assign n4157 = n4148 & n4156;
  assign n4158 = n3408 & n4157;
  assign n4159 = n773 & n4158;
  assign n4160 = n235 & n4159;
  assign n4161 = n454 & n4160;
  assign n4162 = n1040 & n4161;
  assign n4163 = ~n397 & n4162;
  assign n4164 = ~n354 & n4163;
  assign n4165 = ~n1102 & n4164;
  assign n4166 = ~n327 & n4165;
  assign n4167 = ~n403 & n4166;
  assign n4168 = n1524 & n4167;
  assign n4169 = ~n326 & n4168;
  assign n4170 = ~n438 & n4169;
  assign n4171 = ~n201 & n4170;
  assign n4172 = ~n4121 & ~n4171;
  assign n4173 = n4121 & n4171;
  assign n4174 = ~n4172 & ~n4173;
  assign n4175 = ~ a[17]  & n4174;
  assign n4176 = ~n4172 & ~n4175;
  assign n4177 = n3146 & ~n4176;
  assign n4178 = n2916 & ~n2918;
  assign n4179 = ~n2919 & ~n4178;
  assign n4180 = n75 & n4179;
  assign n4181 = ~n710 & n3020;
  assign n4182 = ~n958 & n3023;
  assign n4183 = ~n867 & n3028;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = ~n4181 & n4184;
  assign n4186 = ~n4180 & n4185;
  assign n4187 = ~n3146 & n4176;
  assign n4188 = ~n4177 & ~n4187;
  assign n4189 = ~n4186 & n4188;
  assign n4190 = ~n4177 & ~n4189;
  assign n4191 = ~n4100 & ~n4190;
  assign n4192 = n4100 & n4190;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = ~n4186 & ~n4189;
  assign n4195 = n4188 & ~n4189;
  assign n4196 = ~n4194 & ~n4195;
  assign n4197 = ~ a[17]  & ~n4175;
  assign n4198 = ~n4173 & n4176;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = ~n867 & n3020;
  assign n4201 = ~n958 & n3028;
  assign n4202 = ~n1060 & n3023;
  assign n4203 = n2912 & ~n2914;
  assign n4204 = ~n2915 & ~n4203;
  assign n4205 = n75 & n4204;
  assign n4206 = ~n4202 & ~n4205;
  assign n4207 = ~n4201 & n4206;
  assign n4208 = ~n4200 & n4207;
  assign n4209 = ~n4199 & ~n4208;
  assign n4210 = n2348 & n2515;
  assign n4211 = n977 & n4210;
  assign n4212 = n2090 & n4211;
  assign n4213 = ~n95 & n4212;
  assign n4214 = ~n363 & n4213;
  assign n4215 = ~n449 & n4214;
  assign n4216 = ~n396 & ~n430;
  assign n4217 = ~n236 & ~n1127;
  assign n4218 = ~n875 & n4217;
  assign n4219 = n3085 & n4218;
  assign n4220 = n4216 & n4219;
  assign n4221 = n2132 & n4220;
  assign n4222 = n2301 & n4221;
  assign n4223 = n2202 & n4222;
  assign n4224 = n805 & n4223;
  assign n4225 = n399 & n4224;
  assign n4226 = n227 & n4225;
  assign n4227 = n885 & n4226;
  assign n4228 = ~n136 & n4227;
  assign n4229 = ~n667 & n4228;
  assign n4230 = ~n1102 & n4229;
  assign n4231 = ~n189 & n4230;
  assign n4232 = ~n712 & n4231;
  assign n4233 = ~n496 & n2468;
  assign n4234 = ~n883 & n4233;
  assign n4235 = n3827 & n4234;
  assign n4236 = n778 & n4235;
  assign n4237 = n2017 & n4236;
  assign n4238 = n2740 & n4237;
  assign n4239 = n156 & n4238;
  assign n4240 = ~n123 & n4239;
  assign n4241 = ~n353 & n4240;
  assign n4242 = ~n115 & n4241;
  assign n4243 = ~n233 & n4242;
  assign n4244 = ~n639 & n4243;
  assign n4245 = ~n425 & n4244;
  assign n4246 = ~n99 & n4245;
  assign n4247 = ~n306 & n4246;
  assign n4248 = n541 & n2241;
  assign n4249 = n2330 & n4248;
  assign n4250 = n2507 & n4249;
  assign n4251 = n4247 & n4250;
  assign n4252 = n4232 & n4251;
  assign n4253 = n4215 & n4252;
  assign n4254 = n2635 & n4253;
  assign n4255 = n2682 & n4254;
  assign n4256 = n1781 & n4255;
  assign n4257 = ~n427 & n4256;
  assign n4258 = ~n461 & n4257;
  assign n4259 = ~n228 & n4258;
  assign n4260 = ~n326 & n4259;
  assign n4261 = ~n395 & n4260;
  assign n4262 = ~n714 & n4261;
  assign n4263 = ~n304 & n4262;
  assign n4264 = ~n666 & n4263;
  assign n4265 = ~n886 & n4264;
  assign n4266 = ~n771 & n4265;
  assign n4267 = n4121 & ~n4266;
  assign n4268 = ~n4121 & n4266;
  assign n4269 = ~n150 & ~n155;
  assign n4270 = n250 & n4269;
  assign n4271 = ~n752 & n4270;
  assign n4272 = ~n402 & n4271;
  assign n4273 = ~n430 & n4272;
  assign n4274 = ~n428 & n4273;
  assign n4275 = ~n276 & ~n419;
  assign n4276 = ~n403 & n4275;
  assign n4277 = ~n424 & n4276;
  assign n4278 = ~n170 & n4277;
  assign n4279 = ~n883 & n4278;
  assign n4280 = n1944 & n2684;
  assign n4281 = n4279 & n4280;
  assign n4282 = n4215 & n4281;
  assign n4283 = n4274 & n4282;
  assign n4284 = n1917 & n4283;
  assign n4285 = n773 & n4284;
  assign n4286 = n1237 & n4285;
  assign n4287 = ~n278 & n4286;
  assign n4288 = ~n305 & n4287;
  assign n4289 = ~n146 & n4288;
  assign n4290 = ~n102 & n4289;
  assign n4291 = ~n932 & n4290;
  assign n4292 = ~n200 & n4291;
  assign n4293 = ~n371 & n4292;
  assign n4294 = ~n339 & ~n374;
  assign n4295 = ~n338 & n4294;
  assign n4296 = ~n99 & ~n330;
  assign n4297 = ~n157 & n4296;
  assign n4298 = ~n470 & n4297;
  assign n4299 = n1047 & n2637;
  assign n4300 = n4218 & n4299;
  assign n4301 = n4298 & n4300;
  assign n4302 = n3464 & n4301;
  assign n4303 = n2738 & n4302;
  assign n4304 = n4295 & n4303;
  assign n4305 = ~n123 & n4304;
  assign n4306 = ~n558 & n4305;
  assign n4307 = ~n149 & n4306;
  assign n4308 = ~n527 & n4307;
  assign n4309 = ~n504 & n4308;
  assign n4310 = ~n273 & n4309;
  assign n4311 = ~n564 & n4310;
  assign n4312 = ~n135 & ~n452;
  assign n4313 = ~n283 & n4312;
  assign n4314 = n941 & n4313;
  assign n4315 = n1602 & n4314;
  assign n4316 = ~n154 & n4315;
  assign n4317 = ~n619 & n4316;
  assign n4318 = ~n121 & n4317;
  assign n4319 = ~n594 & n4318;
  assign n4320 = ~n396 & n4319;
  assign n4321 = ~n777 & n4320;
  assign n4322 = ~n326 & n4321;
  assign n4323 = ~n425 & n4322;
  assign n4324 = ~n298 & n4323;
  assign n4325 = ~n791 & n4324;
  assign n4326 = ~n274 & ~n426;
  assign n4327 = ~n633 & n4326;
  assign n4328 = n2371 & n4327;
  assign n4329 = n2073 & n4328;
  assign n4330 = ~n511 & n4329;
  assign n4331 = ~n656 & n4330;
  assign n4332 = ~n657 & n4331;
  assign n4333 = ~n192 & ~n509;
  assign n4334 = ~n340 & n4333;
  assign n4335 = ~n233 & ~n715;
  assign n4336 = n3114 & n4335;
  assign n4337 = n4334 & n4336;
  assign n4338 = n4332 & n4337;
  assign n4339 = n2740 & n4338;
  assign n4340 = n2169 & n4339;
  assign n4341 = n4325 & n4340;
  assign n4342 = n4311 & n4341;
  assign n4343 = n4293 & n4342;
  assign n4344 = n491 & n4343;
  assign n4345 = n1182 & n4344;
  assign n4346 = ~n118 & n4345;
  assign n4347 = ~n689 & n4346;
  assign n4348 = ~n277 & n4347;
  assign n4349 = ~n672 & n4348;
  assign n4350 = ~n86 & n4349;
  assign n4351 = ~n188 & n4350;
  assign n4352 = ~n1246 & n1669;
  assign n4353 = ~n289 & n4352;
  assign n4354 = ~n461 & n4353;
  assign n4355 = ~n363 & n4354;
  assign n4356 = ~n562 & n4355;
  assign n4357 = ~n673 & ~n1306;
  assign n4358 = n1135 & n2334;
  assign n4359 = n4357 & n4358;
  assign n4360 = n1040 & n4359;
  assign n4361 = ~n232 & n4360;
  assign n4362 = ~n255 & n4361;
  assign n4363 = ~n203 & n4362;
  assign n4364 = ~n809 & n4363;
  assign n4365 = ~n239 & n4364;
  assign n4366 = ~n372 & n4365;
  assign n4367 = ~n102 & ~n293;
  assign n4368 = n876 & n2210;
  assign n4369 = n4153 & n4368;
  assign n4370 = n2013 & n4369;
  assign n4371 = n2807 & n4370;
  assign n4372 = n4367 & n4371;
  assign n4373 = ~n169 & n4372;
  assign n4374 = ~n190 & n4373;
  assign n4375 = ~n435 & n4374;
  assign n4376 = n1272 & n4234;
  assign n4377 = n439 & n4376;
  assign n4378 = n4375 & n4377;
  assign n4379 = n3378 & n4378;
  assign n4380 = n1550 & n4379;
  assign n4381 = ~n427 & n4380;
  assign n4382 = ~n420 & n4381;
  assign n4383 = ~n146 & n4382;
  assign n4384 = ~n296 & n4383;
  assign n4385 = ~n980 & n4384;
  assign n4386 = ~n201 & n4385;
  assign n4387 = ~n271 & n4386;
  assign n4388 = ~n249 & n4387;
  assign n4389 = n793 & n3296;
  assign n4390 = n2296 & n4389;
  assign n4391 = n615 & n4390;
  assign n4392 = n1330 & n4391;
  assign n4393 = n827 & n4392;
  assign n4394 = n978 & n4393;
  assign n4395 = n590 & n4394;
  assign n4396 = ~n667 & n4395;
  assign n4397 = ~n355 & n4396;
  assign n4398 = ~n152 & n4397;
  assign n4399 = ~n511 & n4398;
  assign n4400 = ~n594 & n4399;
  assign n4401 = ~n637 & n4400;
  assign n4402 = ~n107 & n4401;
  assign n4403 = ~n601 & n4402;
  assign n4404 = ~n603 & n4403;
  assign n4405 = ~n338 & n4404;
  assign n4406 = n2014 & n3416;
  assign n4407 = n1346 & n4406;
  assign n4408 = n992 & n4407;
  assign n4409 = n1785 & n4408;
  assign n4410 = n4405 & n4409;
  assign n4411 = n4388 & n4410;
  assign n4412 = n4366 & n4411;
  assign n4413 = n4356 & n4412;
  assign n4414 = n774 & n4413;
  assign n4415 = n2698 & n4414;
  assign n4416 = n285 & n4415;
  assign n4417 = ~n236 & n4416;
  assign n4418 = ~n397 & n4417;
  assign n4419 = ~n335 & n4418;
  assign n4420 = ~n563 & n4419;
  assign n4421 = ~n489 & n4420;
  assign n4422 = ~n4351 & ~n4421;
  assign n4423 = n4351 & n4421;
  assign n4424 = ~n4422 & ~n4423;
  assign n4425 = ~ a[14]  & n4424;
  assign n4426 = ~n4422 & ~n4425;
  assign n4427 = n4266 & ~n4426;
  assign n4428 = n2904 & ~n2906;
  assign n4429 = ~n2907 & ~n4428;
  assign n4430 = n75 & n4429;
  assign n4431 = ~n1060 & n3020;
  assign n4432 = ~n1235 & n3023;
  assign n4433 = ~n1178 & n3028;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = ~n4431 & n4434;
  assign n4436 = ~n4430 & n4435;
  assign n4437 = ~n4266 & n4426;
  assign n4438 = ~n4427 & ~n4437;
  assign n4439 = ~n4436 & n4438;
  assign n4440 = ~n4427 & ~n4439;
  assign n4441 = ~n4267 & ~n4440;
  assign n4442 = ~n4268 & n4441;
  assign n4443 = ~n4267 & ~n4442;
  assign n4444 = n4199 & n4208;
  assign n4445 = ~n4209 & ~n4444;
  assign n4446 = ~n4443 & n4445;
  assign n4447 = ~n4209 & ~n4446;
  assign n4448 = ~n4196 & ~n4447;
  assign n4449 = n4196 & n4447;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = ~n3012 & n3457;
  assign n4452 = ~n587 & n3542;
  assign n4453 = ~n392 & n3606;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = ~n4451 & n4454;
  assign n4456 = ~n3368 & n4455;
  assign n4457 = ~n3018 & n4455;
  assign n4458 = ~n4456 & ~n4457;
  assign n4459 =  a[29]  & ~n4458;
  assign n4460 = ~ a[29]  & n4458;
  assign n4461 = ~n4459 & ~n4460;
  assign n4462 = n4450 & ~n4461;
  assign n4463 = ~n4448 & ~n4462;
  assign n4464 = n4193 & ~n4463;
  assign n4465 = ~n4191 & ~n4464;
  assign n4466 = ~n4097 & ~n4465;
  assign n4467 = ~n4094 & ~n4466;
  assign n4468 = ~n3361 & n3632;
  assign n4469 = ~n3633 & ~n4468;
  assign n4470 = ~n4467 & n4469;
  assign n4471 = n3884 & ~n4045;
  assign n4472 = ~n3805 & n3967;
  assign n4473 = ~n3964 & n4046;
  assign n4474 = ~n4472 & ~n4473;
  assign n4475 = ~n4471 & n4474;
  assign n4476 = n4057 & ~n4059;
  assign n4477 = ~n4060 & ~n4476;
  assign n4478 = n4050 & n4477;
  assign n4479 = n4475 & ~n4478;
  assign n4480 =  a[26]  & ~n4479;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 =  a[26]  & ~n4480;
  assign n4483 = ~n4481 & ~n4482;
  assign n4484 = ~n4467 & ~n4470;
  assign n4485 = n4469 & ~n4470;
  assign n4486 = ~n4484 & ~n4485;
  assign n4487 = ~n4483 & ~n4486;
  assign n4488 = ~n4470 & ~n4487;
  assign n4489 = ~n714 & n2014;
  assign n4490 = ~n243 & n4489;
  assign n4491 = ~n145 & n4490;
  assign n4492 = ~n466 & n4491;
  assign n4493 = ~n205 & n4492;
  assign n4494 = n1388 & n1785;
  assign n4495 = n604 & n4494;
  assign n4496 = n2170 & n4495;
  assign n4497 = ~n173 & n4496;
  assign n4498 = ~n144 & n4497;
  assign n4499 = ~n394 & n4498;
  assign n4500 = ~n306 & n4499;
  assign n4501 = ~n157 & n4500;
  assign n4502 = ~n375 & n4501;
  assign n4503 = n133 & n4502;
  assign n4504 = n4493 & n4503;
  assign n4505 = n2346 & n4504;
  assign n4506 = n1046 & n4505;
  assign n4507 = n1761 & n4506;
  assign n4508 = n1367 & n4507;
  assign n4509 = ~n274 & n4508;
  assign n4510 = ~n589 & n4509;
  assign n4511 = ~n468 & n4510;
  assign n4512 = n3972 & n4511;
  assign n4513 = ~n296 & n4512;
  assign n4514 = ~n601 & n4513;
  assign n4515 = n3839 & n4514;
  assign n4516 = ~n4062 & ~n4065;
  assign n4517 = ~n3877 & ~n4515;
  assign n4518 = n3877 & n4515;
  assign n4519 = ~n4517 & ~n4518;
  assign n4520 = ~n4516 & n4519;
  assign n4521 = n3877 & ~n4520;
  assign n4522 = ~n4515 & ~n4521;
  assign n4523 = ~ a[21]  &  a[22] ;
  assign n4524 =  a[21]  & ~ a[22] ;
  assign n4525 = ~n4523 & ~n4524;
  assign n4526 =  a[20]  & ~ a[21] ;
  assign n4527 = ~ a[20]  &  a[21] ;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = ~ a[22]  &  a[23] ;
  assign n4530 =  a[22]  & ~ a[23] ;
  assign n4531 = ~n4529 & ~n4530;
  assign n4532 = n4528 & ~n4531;
  assign n4533 = n4525 & n4532;
  assign n4534 = ~n4515 & n4533;
  assign n4535 = ~n4522 & ~n4534;
  assign n4536 = ~n4528 & ~n4531;
  assign n4537 = ~n4534 & ~n4536;
  assign n4538 = ~n4535 & ~n4537;
  assign n4539 =  a[23]  & ~n4538;
  assign n4540 = ~ a[23]  & n4538;
  assign n4541 = ~n4539 & ~n4540;
  assign n4542 = ~n4488 & ~n4541;
  assign n4543 = n4488 & n4541;
  assign n4544 = ~n4542 & ~n4543;
  assign n4545 = ~n4077 & n4544;
  assign n4546 = ~n4077 & ~n4545;
  assign n4547 = n4544 & ~n4545;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = n4097 & n4465;
  assign n4550 = ~n4466 & ~n4549;
  assign n4551 = n3884 & ~n3964;
  assign n4552 = ~n3456 & n3967;
  assign n4553 = ~n3805 & n4046;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = ~n4551 & n4554;
  assign n4556 = ~n4050 & n4555;
  assign n4557 = n4053 & ~n4055;
  assign n4558 = ~n4056 & ~n4557;
  assign n4559 = n4555 & ~n4558;
  assign n4560 = ~n4556 & ~n4559;
  assign n4561 =  a[26]  & ~n4560;
  assign n4562 = ~ a[26]  & n4560;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = n4550 & ~n4563;
  assign n4565 = ~n3805 & n3884;
  assign n4566 = ~n3605 & n3967;
  assign n4567 = ~n3456 & n4046;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = ~n4565 & n4568;
  assign n4570 = n3818 & n4050;
  assign n4571 = n4569 & ~n4570;
  assign n4572 =  a[26]  & ~n4571;
  assign n4573 =  a[26]  & ~n4572;
  assign n4574 = ~n4571 & ~n4572;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = ~n4193 & n4463;
  assign n4577 = ~n4464 & ~n4576;
  assign n4578 = n3457 & ~n3539;
  assign n4579 = ~n392 & n3542;
  assign n4580 = ~n3012 & n3606;
  assign n4581 = ~n4579 & ~n4580;
  assign n4582 = ~n4578 & n4581;
  assign n4583 = ~n3368 & n4582;
  assign n4584 = ~n3715 & n4582;
  assign n4585 = ~n4583 & ~n4584;
  assign n4586 =  a[29]  & ~n4585;
  assign n4587 = ~ a[29]  & n4585;
  assign n4588 = ~n4586 & ~n4587;
  assign n4589 = n4577 & ~n4588;
  assign n4590 = ~n4577 & n4588;
  assign n4591 = ~n4589 & ~n4590;
  assign n4592 = ~n4575 & n4591;
  assign n4593 = ~n4589 & ~n4592;
  assign n4594 = n4550 & ~n4564;
  assign n4595 = ~n4563 & ~n4564;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = ~n4593 & ~n4596;
  assign n4598 = ~n4564 & ~n4597;
  assign n4599 = n4483 & ~n4485;
  assign n4600 = ~n4484 & n4599;
  assign n4601 = ~n4487 & ~n4600;
  assign n4602 = ~n4598 & n4601;
  assign n4603 = ~n3877 & n4533;
  assign n4604 = ~n4525 & n4528;
  assign n4605 = ~n4515 & n4604;
  assign n4606 = ~n4603 & ~n4605;
  assign n4607 = ~n4517 & ~n4520;
  assign n4608 = n4515 & n4607;
  assign n4609 = ~n4522 & ~n4608;
  assign n4610 = n4536 & n4609;
  assign n4611 = n4606 & ~n4610;
  assign n4612 =  a[23]  & ~n4611;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 =  a[23]  & ~n4612;
  assign n4615 = ~n4613 & ~n4614;
  assign n4616 = n4598 & ~n4601;
  assign n4617 = ~n4602 & ~n4616;
  assign n4618 = ~n4615 & n4617;
  assign n4619 = ~n4602 & ~n4618;
  assign n4620 = n4548 & n4619;
  assign n4621 = ~n4548 & ~n4619;
  assign n4622 = ~n4620 & ~n4621;
  assign n4623 = n4591 & ~n4592;
  assign n4624 = ~n4575 & ~n4592;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~n4440 & ~n4442;
  assign n4627 = ~n4268 & n4443;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = ~n958 & n3020;
  assign n4630 = ~n1060 & n3028;
  assign n4631 = ~n1178 & n3023;
  assign n4632 = n2908 & ~n2910;
  assign n4633 = ~n2911 & ~n4632;
  assign n4634 = n75 & n4633;
  assign n4635 = ~n4631 & ~n4634;
  assign n4636 = ~n4630 & n4635;
  assign n4637 = ~n4629 & n4636;
  assign n4638 = ~n4628 & ~n4637;
  assign n4639 = ~n587 & n3457;
  assign n4640 = ~n867 & n3542;
  assign n4641 = ~n710 & n3606;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = ~n4639 & n4642;
  assign n4644 = n3331 & n3368;
  assign n4645 = n4643 & ~n4644;
  assign n4646 =  a[29]  & ~n4645;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 =  a[29]  & ~n4646;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = ~n4628 & ~n4638;
  assign n4651 = ~n4637 & ~n4638;
  assign n4652 = ~n4650 & ~n4651;
  assign n4653 = ~n4649 & ~n4652;
  assign n4654 = ~n4638 & ~n4653;
  assign n4655 = n4443 & ~n4445;
  assign n4656 = ~n4446 & ~n4655;
  assign n4657 = ~n4654 & n4656;
  assign n4658 = ~n392 & n3457;
  assign n4659 = ~n710 & n3542;
  assign n4660 = ~n587 & n3606;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = ~n4658 & n4661;
  assign n4663 = n3347 & n3368;
  assign n4664 = n4662 & ~n4663;
  assign n4665 =  a[29]  & ~n4664;
  assign n4666 =  a[29]  & ~n4665;
  assign n4667 = ~n4664 & ~n4665;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = n4654 & ~n4656;
  assign n4670 = ~n4657 & ~n4669;
  assign n4671 = ~n4668 & n4670;
  assign n4672 = ~n4657 & ~n4671;
  assign n4673 = ~n4450 & n4461;
  assign n4674 = ~n4462 & ~n4673;
  assign n4675 = ~n4672 & n4674;
  assign n4676 = n4672 & ~n4674;
  assign n4677 = ~n4675 & ~n4676;
  assign n4678 = ~n3456 & n3884;
  assign n4679 = ~n3539 & n3967;
  assign n4680 = ~n3605 & n4046;
  assign n4681 = ~n4679 & ~n4680;
  assign n4682 = ~n4678 & n4681;
  assign n4683 = n3627 & n4050;
  assign n4684 = n4682 & ~n4683;
  assign n4685 =  a[26]  & ~n4684;
  assign n4686 =  a[26]  & ~n4685;
  assign n4687 = ~n4684 & ~n4685;
  assign n4688 = ~n4686 & ~n4687;
  assign n4689 = n4677 & ~n4688;
  assign n4690 = ~n4675 & ~n4689;
  assign n4691 = ~n4625 & ~n4690;
  assign n4692 = n4625 & n4690;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = ~n4528 & n4531;
  assign n4695 = ~n3877 & n4694;
  assign n4696 = ~n3964 & n4533;
  assign n4697 = ~n4045 & n4604;
  assign n4698 = ~n4696 & ~n4697;
  assign n4699 = ~n4695 & n4698;
  assign n4700 = n4067 & n4536;
  assign n4701 = n4699 & ~n4700;
  assign n4702 =  a[23]  & ~n4701;
  assign n4703 =  a[23]  & ~n4702;
  assign n4704 = ~n4701 & ~n4702;
  assign n4705 = ~n4703 & ~n4704;
  assign n4706 = n4693 & ~n4705;
  assign n4707 = ~n4691 & ~n4706;
  assign n4708 = ~n4515 & n4694;
  assign n4709 = ~n4045 & n4533;
  assign n4710 = ~n3877 & n4604;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = ~n4708 & n4711;
  assign n4713 = ~n4536 & n4712;
  assign n4714 = n4516 & ~n4519;
  assign n4715 = ~n4520 & ~n4714;
  assign n4716 = n4712 & ~n4715;
  assign n4717 = ~n4713 & ~n4716;
  assign n4718 =  a[23]  & ~n4717;
  assign n4719 = ~ a[23]  & n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~n4707 & ~n4720;
  assign n4722 = n4707 & n4720;
  assign n4723 = ~n4721 & ~n4722;
  assign n4724 = ~n4593 & ~n4597;
  assign n4725 = ~n4596 & ~n4597;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = n4723 & ~n4726;
  assign n4728 = ~n4721 & ~n4727;
  assign n4729 = n4615 & ~n4617;
  assign n4730 = ~n4618 & ~n4729;
  assign n4731 = ~n4728 & n4730;
  assign n4732 = n4723 & ~n4727;
  assign n4733 = ~n4726 & ~n4727;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = n4677 & ~n4689;
  assign n4736 = ~n4688 & ~n4689;
  assign n4737 = ~n4735 & ~n4736;
  assign n4738 = n4670 & ~n4671;
  assign n4739 = ~n4668 & ~n4671;
  assign n4740 = ~n4738 & ~n4739;
  assign n4741 = ~n3605 & n3884;
  assign n4742 = ~n3012 & n3967;
  assign n4743 = ~n3539 & n4046;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = ~n4741 & n4744;
  assign n4746 = ~n4050 & n4745;
  assign n4747 = ~n4084 & n4745;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 =  a[26]  & ~n4748;
  assign n4750 = ~ a[26]  & n4748;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~n4740 & ~n4751;
  assign n4753 = ~n4649 & ~n4653;
  assign n4754 = ~n4652 & ~n4653;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = ~n4436 & ~n4439;
  assign n4757 = n4438 & ~n4439;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~ a[14]  & ~n4425;
  assign n4760 = ~n4423 & n4426;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = ~n617 & n3043;
  assign n4763 = ~n154 & n4762;
  assign n4764 = ~n641 & n4763;
  assign n4765 = ~n328 & n4764;
  assign n4766 = ~n394 & n4765;
  assign n4767 = ~n666 & n4766;
  assign n4768 = ~n564 & n3490;
  assign n4769 = ~n886 & n4768;
  assign n4770 = n333 & n1389;
  assign n4771 = ~n449 & n4770;
  assign n4772 = n2361 & n4771;
  assign n4773 = n4769 & n4772;
  assign n4774 = n141 & n4773;
  assign n4775 = n1181 & n4774;
  assign n4776 = n874 & n4775;
  assign n4777 = n968 & n4776;
  assign n4778 = n3252 & n4777;
  assign n4779 = n1827 & n4778;
  assign n4780 = n2583 & n4779;
  assign n4781 = n4101 & n4780;
  assign n4782 = ~n169 & n4781;
  assign n4783 = ~n286 & n4782;
  assign n4784 = ~n589 & n4783;
  assign n4785 = ~n252 & n4784;
  assign n4786 = ~n335 & ~n367;
  assign n4787 = ~n375 & ~n511;
  assign n4788 = ~n304 & n4787;
  assign n4789 = n2154 & n4788;
  assign n4790 = ~n1306 & n4789;
  assign n4791 = ~n397 & n4790;
  assign n4792 = ~n189 & n4791;
  assign n4793 = ~n233 & n4792;
  assign n4794 = ~n161 & n4793;
  assign n4795 = ~n205 & ~n275;
  assign n4796 = ~n961 & n4795;
  assign n4797 = ~n249 & n4796;
  assign n4798 = n1761 & n4367;
  assign n4799 = ~n715 & n4798;
  assign n4800 = n4797 & n4799;
  assign n4801 = n297 & n4800;
  assign n4802 = n439 & n4801;
  assign n4803 = n4794 & n4802;
  assign n4804 = n4786 & n4803;
  assign n4805 = n933 & n4804;
  assign n4806 = n2219 & n4805;
  assign n4807 = n341 & n4806;
  assign n4808 = ~n469 & n4807;
  assign n4809 = ~n276 & n4808;
  assign n4810 = ~n557 & n4809;
  assign n4811 = ~n602 & n4810;
  assign n4812 = ~n150 & n4811;
  assign n4813 = ~n416 & n4812;
  assign n4814 = ~n191 & n4813;
  assign n4815 = ~n791 & n4814;
  assign n4816 = ~n164 & ~n558;
  assign n4817 = ~n537 & n4816;
  assign n4818 = ~n200 & n4817;
  assign n4819 = ~n672 & n4818;
  assign n4820 = n2584 & n2721;
  assign n4821 = n4819 & n4820;
  assign n4822 = n1726 & n4821;
  assign n4823 = n570 & n4822;
  assign n4824 = ~n1011 & n4823;
  assign n4825 = ~n290 & n4824;
  assign n4826 = ~n246 & n4825;
  assign n4827 = ~n393 & n4826;
  assign n4828 = ~n496 & ~n884;
  assign n4829 = n1973 & n4828;
  assign n4830 = n4827 & n4829;
  assign n4831 = n4815 & n4830;
  assign n4832 = n1928 & n4831;
  assign n4833 = n4785 & n4832;
  assign n4834 = n4767 & n4833;
  assign n4835 = n1576 & n4834;
  assign n4836 = n423 & n4835;
  assign n4837 = n2467 & n4836;
  assign n4838 = ~n667 & n4837;
  assign n4839 = ~n91 & n4838;
  assign n4840 = ~n243 & n4839;
  assign n4841 = ~n536 & n4840;
  assign n4842 = ~n283 & n4841;
  assign n4843 = ~n237 & n4842;
  assign n4844 = ~n271 & n4843;
  assign n4845 = n4351 & ~n4844;
  assign n4846 = ~n4351 & n4844;
  assign n4847 = n2896 & ~n2898;
  assign n4848 = ~n2899 & ~n4847;
  assign n4849 = n75 & n4848;
  assign n4850 = ~n1235 & n3020;
  assign n4851 = ~n1472 & n3023;
  assign n4852 = ~n1364 & n3028;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~n4850 & n4853;
  assign n4855 = ~n4849 & n4854;
  assign n4856 = ~n4845 & ~n4855;
  assign n4857 = ~n4846 & n4856;
  assign n4858 = ~n4845 & ~n4857;
  assign n4859 = ~n4761 & ~n4858;
  assign n4860 = n2900 & ~n2902;
  assign n4861 = ~n2903 & ~n4860;
  assign n4862 = n75 & n4861;
  assign n4863 = ~n1178 & n3020;
  assign n4864 = ~n1364 & n3023;
  assign n4865 = ~n1235 & n3028;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = ~n4863 & n4866;
  assign n4868 = ~n4862 & n4867;
  assign n4869 = n4761 & n4858;
  assign n4870 = ~n4859 & ~n4869;
  assign n4871 = ~n4868 & n4870;
  assign n4872 = ~n4859 & ~n4871;
  assign n4873 = ~n4758 & ~n4872;
  assign n4874 = n4758 & n4872;
  assign n4875 = ~n4873 & ~n4874;
  assign n4876 = ~n710 & n3457;
  assign n4877 = ~n958 & n3542;
  assign n4878 = ~n867 & n3606;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~n4876 & n4879;
  assign n4881 = ~n3368 & n4880;
  assign n4882 = ~n4179 & n4880;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 =  a[29]  & ~n4883;
  assign n4885 = ~ a[29]  & n4883;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = n4875 & ~n4886;
  assign n4888 = ~n4873 & ~n4887;
  assign n4889 = ~n4755 & ~n4888;
  assign n4890 = n4755 & n4888;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = ~n3539 & n3884;
  assign n4893 = ~n392 & n3967;
  assign n4894 = ~n3012 & n4046;
  assign n4895 = ~n4893 & ~n4894;
  assign n4896 = ~n4892 & n4895;
  assign n4897 = n3715 & n4050;
  assign n4898 = n4896 & ~n4897;
  assign n4899 =  a[26]  & ~n4898;
  assign n4900 =  a[26]  & ~n4899;
  assign n4901 = ~n4898 & ~n4899;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = n4891 & ~n4902;
  assign n4904 = ~n4889 & ~n4903;
  assign n4905 = n4740 & n4751;
  assign n4906 = ~n4752 & ~n4905;
  assign n4907 = ~n4904 & n4906;
  assign n4908 = ~n4752 & ~n4907;
  assign n4909 = ~n4737 & ~n4908;
  assign n4910 = n4737 & n4908;
  assign n4911 = ~n4909 & ~n4910;
  assign n4912 = ~n4045 & n4694;
  assign n4913 = ~n3805 & n4533;
  assign n4914 = ~n3964 & n4604;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = ~n4912 & n4915;
  assign n4917 = n4477 & n4536;
  assign n4918 = n4916 & ~n4917;
  assign n4919 =  a[23]  & ~n4918;
  assign n4920 =  a[23]  & ~n4919;
  assign n4921 = ~n4918 & ~n4919;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = n4911 & ~n4922;
  assign n4924 = ~n4909 & ~n4923;
  assign n4925 = ~ a[18]  &  a[19] ;
  assign n4926 =  a[18]  & ~ a[19] ;
  assign n4927 = ~n4925 & ~n4926;
  assign n4928 =  a[19]  & ~ a[20] ;
  assign n4929 = ~ a[19]  &  a[20] ;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 =  a[17]  & ~ a[18] ;
  assign n4932 = ~ a[17]  &  a[18] ;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = ~n4930 & n4933;
  assign n4935 = n4927 & n4934;
  assign n4936 = ~n4515 & n4935;
  assign n4937 = ~n4522 & ~n4936;
  assign n4938 = ~n4930 & ~n4933;
  assign n4939 = ~n4936 & ~n4938;
  assign n4940 = ~n4937 & ~n4939;
  assign n4941 =  a[20]  & ~n4940;
  assign n4942 = ~ a[20]  & n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4924 & ~n4943;
  assign n4945 = n4693 & ~n4706;
  assign n4946 = ~n4705 & ~n4706;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = n4924 & n4943;
  assign n4949 = ~n4944 & ~n4948;
  assign n4950 = ~n4947 & n4949;
  assign n4951 = ~n4944 & ~n4950;
  assign n4952 = ~n4734 & ~n4951;
  assign n4953 = n4734 & n4951;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = ~n4947 & ~n4950;
  assign n4956 = n4949 & ~n4950;
  assign n4957 = ~n4955 & ~n4956;
  assign n4958 = n4911 & ~n4923;
  assign n4959 = ~n4922 & ~n4923;
  assign n4960 = ~n4958 & ~n4959;
  assign n4961 = ~n3964 & n4694;
  assign n4962 = ~n3456 & n4533;
  assign n4963 = ~n3805 & n4604;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = ~n4961 & n4964;
  assign n4966 = n4536 & n4558;
  assign n4967 = n4965 & ~n4966;
  assign n4968 =  a[23]  & ~n4967;
  assign n4969 = ~n4967 & ~n4968;
  assign n4970 =  a[23]  & ~n4968;
  assign n4971 = ~n4969 & ~n4970;
  assign n4972 = n4904 & ~n4906;
  assign n4973 = ~n4907 & ~n4972;
  assign n4974 = ~n4971 & n4973;
  assign n4975 = ~n4971 & ~n4974;
  assign n4976 = n4973 & ~n4974;
  assign n4977 = ~n4975 & ~n4976;
  assign n4978 = n4891 & ~n4903;
  assign n4979 = ~n4902 & ~n4903;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = ~n867 & n3457;
  assign n4982 = ~n1060 & n3542;
  assign n4983 = ~n958 & n3606;
  assign n4984 = ~n4982 & ~n4983;
  assign n4985 = ~n4981 & n4984;
  assign n4986 = n3368 & n4204;
  assign n4987 = n4985 & ~n4986;
  assign n4988 =  a[29]  & ~n4987;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 =  a[29]  & ~n4988;
  assign n4991 = ~n4989 & ~n4990;
  assign n4992 = ~n4868 & ~n4871;
  assign n4993 = n4870 & ~n4871;
  assign n4994 = ~n4992 & ~n4993;
  assign n4995 = ~n4991 & ~n4994;
  assign n4996 = ~n4991 & ~n4995;
  assign n4997 = ~n4994 & ~n4995;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = ~n4855 & ~n4857;
  assign n5000 = ~n4846 & n4858;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = ~n394 & ~n1062;
  assign n5003 = n2546 & n5002;
  assign n5004 = n4357 & n5003;
  assign n5005 = n3438 & n5004;
  assign n5006 = n3886 & n5005;
  assign n5007 = n421 & n5006;
  assign n5008 = n1237 & n5007;
  assign n5009 = ~n305 & n5008;
  assign n5010 = ~n302 & n5009;
  assign n5011 = ~n589 & n5010;
  assign n5012 = ~n468 & n5011;
  assign n5013 = ~n883 & n5012;
  assign n5014 = ~n364 & n1709;
  assign n5015 = ~n121 & n5014;
  assign n5016 = ~n422 & n5015;
  assign n5017 = ~n130 & n5016;
  assign n5018 = ~n325 & n5017;
  assign n5019 = ~n158 & n5018;
  assign n5020 = ~n170 & ~n825;
  assign n5021 = ~n519 & n5020;
  assign n5022 = n1331 & n1861;
  assign n5023 = n5021 & n5022;
  assign n5024 = n811 & n5023;
  assign n5025 = n5019 & n5024;
  assign n5026 = n3163 & n5025;
  assign n5027 = ~n154 & n5026;
  assign n5028 = ~n135 & n5027;
  assign n5029 = ~n1102 & n5028;
  assign n5030 = ~n402 & n5029;
  assign n5031 = ~n290 & n5030;
  assign n5032 = ~n374 & n5031;
  assign n5033 = ~n689 & n5032;
  assign n5034 = ~n231 & n5033;
  assign n5035 = ~n304 & ~n513;
  assign n5036 = ~n251 & n5035;
  assign n5037 = ~n339 & ~n398;
  assign n5038 = ~n283 & n5037;
  assign n5039 = n979 & n2406;
  assign n5040 = ~n1072 & n5039;
  assign n5041 = n812 & n5040;
  assign n5042 = n5038 & n5041;
  assign n5043 = n5036 & n5042;
  assign n5044 = n4216 & n5043;
  assign n5045 = n4332 & n5044;
  assign n5046 = n1610 & n5045;
  assign n5047 = n2979 & n5046;
  assign n5048 = n5034 & n5047;
  assign n5049 = n5013 & n5048;
  assign n5050 = ~n752 & n5049;
  assign n5051 = ~n1101 & n5050;
  assign n5052 = ~n201 & n5051;
  assign n5053 = ~n562 & n5052;
  assign n5054 = ~n511 & ~n746;
  assign n5055 = ~n283 & n5054;
  assign n5056 = ~n562 & n5055;
  assign n5057 = n2608 & n3043;
  assign n5058 = n5056 & n5057;
  assign n5059 = n621 & n5058;
  assign n5060 = n896 & n5059;
  assign n5061 = ~n403 & n5060;
  assign n5062 = ~n416 & n5061;
  assign n5063 = ~n144 & n5062;
  assign n5064 = ~n225 & ~n716;
  assign n5065 = ~n280 & ~n847;
  assign n5066 = ~n402 & n5065;
  assign n5067 = n5064 & n5066;
  assign n5068 = n1249 & n5067;
  assign n5069 = n5063 & n5068;
  assign n5070 = n664 & n5069;
  assign n5071 = n1668 & n5070;
  assign n5072 = n1667 & n5071;
  assign n5073 = n356 & n5072;
  assign n5074 = n1040 & n5073;
  assign n5075 = ~n617 & n5074;
  assign n5076 = ~n169 & n5075;
  assign n5077 = ~n329 & n5076;
  assign n5078 = ~n335 & n5077;
  assign n5079 = ~n803 & n5078;
  assign n5080 = ~n1203 & n5079;
  assign n5081 = ~n375 & n5080;
  assign n5082 = ~n158 & n5081;
  assign n5083 = ~n298 & ~n825;
  assign n5084 = ~n130 & n5083;
  assign n5085 = ~n493 & n5084;
  assign n5086 = n1012 & n1107;
  assign n5087 = n3663 & n5086;
  assign n5088 = n789 & n5087;
  assign n5089 = n811 & n5088;
  assign n5090 = n3094 & n5089;
  assign n5091 = n5085 & n5090;
  assign n5092 = n2170 & n5091;
  assign n5093 = n5082 & n5092;
  assign n5094 = n5013 & n5093;
  assign n5095 = n508 & n5094;
  assign n5096 = n116 & n5095;
  assign n5097 = n418 & n5096;
  assign n5098 = ~n278 & n5097;
  assign n5099 = ~n506 & n5098;
  assign n5100 = ~n594 & n5099;
  assign n5101 = ~n286 & n5100;
  assign n5102 = ~n424 & n5101;
  assign n5103 = ~n932 & n5102;
  assign n5104 = ~n340 & n5103;
  assign n5105 = ~n337 & n5104;
  assign n5106 = ~n429 & n5105;
  assign n5107 = ~n5053 & ~n5106;
  assign n5108 = n5053 & n5106;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = ~ a[11]  & n5109;
  assign n5111 = ~n5107 & ~n5110;
  assign n5112 = n4351 & ~n5111;
  assign n5113 = n2892 & ~n2894;
  assign n5114 = ~n2895 & ~n5113;
  assign n5115 = n75 & n5114;
  assign n5116 = ~n1364 & n3020;
  assign n5117 = ~n1572 & n3023;
  assign n5118 = ~n1472 & n3028;
  assign n5119 = ~n5117 & ~n5118;
  assign n5120 = ~n5116 & n5119;
  assign n5121 = ~n5115 & n5120;
  assign n5122 = ~n4351 & n5111;
  assign n5123 = ~n5112 & ~n5122;
  assign n5124 = ~n5121 & n5123;
  assign n5125 = ~n5112 & ~n5124;
  assign n5126 = ~n5001 & ~n5125;
  assign n5127 = n5001 & n5125;
  assign n5128 = ~n5126 & ~n5127;
  assign n5129 = ~n5121 & ~n5124;
  assign n5130 = n5123 & ~n5124;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = ~ a[11]  & ~n5110;
  assign n5133 = ~n5108 & n5111;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = ~n1472 & n3020;
  assign n5136 = ~n1572 & n3028;
  assign n5137 = ~n1665 & n3023;
  assign n5138 = n2888 & ~n2890;
  assign n5139 = ~n2891 & ~n5138;
  assign n5140 = n75 & n5139;
  assign n5141 = ~n5137 & ~n5140;
  assign n5142 = ~n5136 & n5141;
  assign n5143 = ~n5135 & n5142;
  assign n5144 = ~n5134 & ~n5143;
  assign n5145 = ~n115 & n1183;
  assign n5146 = ~n107 & n5145;
  assign n5147 = ~n205 & n5146;
  assign n5148 = ~n564 & n5147;
  assign n5149 = ~n428 & n1523;
  assign n5150 = ~n270 & n5149;
  assign n5151 = ~n168 & n1330;
  assign n5152 = ~n252 & n5151;
  assign n5153 = n5150 & n5152;
  assign n5154 = n921 & n5153;
  assign n5155 = n5148 & n5154;
  assign n5156 = n1635 & n5155;
  assign n5157 = n3651 & n5156;
  assign n5158 = n1585 & n5157;
  assign n5159 = n1915 & n5158;
  assign n5160 = n2484 & n5159;
  assign n5161 = n770 & n5160;
  assign n5162 = ~n1072 & n5161;
  assign n5163 = ~n514 & n5162;
  assign n5164 = ~n290 & n5163;
  assign n5165 = ~n825 & n5164;
  assign n5166 = ~n673 & n5165;
  assign n5167 = ~n537 & n5166;
  assign n5168 = ~n325 & n5167;
  assign n5169 = n5053 & ~n5168;
  assign n5170 = ~n5053 & n5168;
  assign n5171 = ~n713 & ~n1101;
  assign n5172 = ~n328 & n1128;
  assign n5173 = ~n287 & n5172;
  assign n5174 = n2278 & n5173;
  assign n5175 = n897 & n5174;
  assign n5176 = n4356 & n5175;
  assign n5177 = n512 & n5176;
  assign n5178 = n654 & n5177;
  assign n5179 = n356 & n5178;
  assign n5180 = n3163 & n5179;
  assign n5181 = ~n571 & n5180;
  assign n5182 = ~n396 & n5181;
  assign n5183 = ~n226 & n5182;
  assign n5184 = ~n639 & n5183;
  assign n5185 = ~n980 & n5184;
  assign n5186 = ~n200 & n5185;
  assign n5187 = ~n272 & n5186;
  assign n5188 = ~n295 & n5187;
  assign n5189 = ~n169 & ~n462;
  assign n5190 = ~n286 & n5189;
  assign n5191 = n2423 & n5190;
  assign n5192 = ~n1011 & n5191;
  assign n5193 = ~n327 & n5192;
  assign n5194 = ~n326 & n2240;
  assign n5195 = ~n673 & n5194;
  assign n5196 = ~n961 & n5195;
  assign n5197 = ~n603 & n5196;
  assign n5198 = ~n366 & n5197;
  assign n5199 = ~n886 & n5198;
  assign n5200 = ~n175 & ~n453;
  assign n5201 = ~n449 & n5200;
  assign n5202 = ~n236 & n5201;
  assign n5203 = ~n746 & n5202;
  assign n5204 = ~n229 & n5203;
  assign n5205 = ~n150 & n5204;
  assign n5206 = ~n438 & n5205;
  assign n5207 = ~n243 & n5206;
  assign n5208 = ~n372 & n5207;
  assign n5209 = ~n655 & n5208;
  assign n5210 = n2297 & n4313;
  assign n5211 = n593 & n5210;
  assign n5212 = n1024 & n5211;
  assign n5213 = n1131 & n5212;
  assign n5214 = n5209 & n5213;
  assign n5215 = n5199 & n5214;
  assign n5216 = ~n111 & n5215;
  assign n5217 = ~n620 & n5216;
  assign n5218 = ~n417 & n5217;
  assign n5219 = ~n167 & n5218;
  assign n5220 = ~n173 & n5219;
  assign n5221 = ~n623 & n5220;
  assign n5222 = ~n1104 & n5221;
  assign n5223 = ~n474 & n5222;
  assign n5224 = ~n569 & n5223;
  assign n5225 = n1085 & n2752;
  assign n5226 = n1155 & n5225;
  assign n5227 = n1367 & n5226;
  assign n5228 = ~n330 & n5227;
  assign n5229 = ~n298 & n5228;
  assign n5230 = ~n130 & n5229;
  assign n5231 = ~n712 & n5230;
  assign n5232 = ~n532 & n5231;
  assign n5233 = ~n81 & n5232;
  assign n5234 = n1732 & n2133;
  assign n5235 = ~n232 & n5234;
  assign n5236 = ~n255 & n5235;
  assign n5237 = ~n299 & n5236;
  assign n5238 = ~n527 & n5237;
  assign n5239 = ~n158 & n5238;
  assign n5240 = n636 & n5066;
  assign n5241 = n1819 & n5240;
  assign n5242 = n5239 & n5241;
  assign n5243 = n5233 & n5242;
  assign n5244 = n5224 & n5243;
  assign n5245 = n5193 & n5244;
  assign n5246 = n5188 & n5245;
  assign n5247 = ~n602 & n5246;
  assign n5248 = n5171 & n5247;
  assign n5249 = ~n339 & n5248;
  assign n5250 = ~n145 & n5249;
  assign n5251 = ~n201 & n5250;
  assign n5252 = ~n666 & n5251;
  assign n5253 = ~n337 & n5252;
  assign n5254 = ~n429 & n5253;
  assign n5255 = n2424 & n3040;
  assign n5256 = n2021 & n5255;
  assign n5257 = ~n364 & n5256;
  assign n5258 = ~n355 & n5257;
  assign n5259 = ~n152 & n5258;
  assign n5260 = ~n115 & n5259;
  assign n5261 = ~n884 & n5260;
  assign n5262 = ~n191 & n5261;
  assign n5263 = ~n1104 & n5262;
  assign n5264 = ~n449 & n5263;
  assign n5265 = n634 & n937;
  assign n5266 = ~n275 & n5265;
  assign n5267 = ~n240 & n5266;
  assign n5268 = ~n188 & n5267;
  assign n5269 = ~n249 & n5268;
  assign n5270 = n202 & ~n513;
  assign n5271 = ~n428 & n5270;
  assign n5272 = n3268 & n5271;
  assign n5273 = n593 & n5272;
  assign n5274 = n5269 & n5273;
  assign n5275 = n5264 & n5274;
  assign n5276 = n873 & n5275;
  assign n5277 = n872 & n5276;
  assign n5278 = n2346 & n5277;
  assign n5279 = n1575 & n5278;
  assign n5280 = n621 & n5279;
  assign n5281 = ~n1306 & n5280;
  assign n5282 = ~n284 & n5281;
  assign n5283 = ~n425 & n5282;
  assign n5284 = ~n306 & n5283;
  assign n5285 = ~n157 & n5284;
  assign n5286 = ~n519 & n5285;
  assign n5287 = n1604 & n2508;
  assign n5288 = n1103 & n5287;
  assign n5289 = n665 & n5288;
  assign n5290 = ~n123 & n5289;
  assign n5291 = ~n107 & n5290;
  assign n5292 = ~n305 & n5291;
  assign n5293 = ~n287 & n5292;
  assign n5294 = ~n490 & n5293;
  assign n5295 = ~n375 & n5294;
  assign n5296 = ~n277 & n5295;
  assign n5297 = ~n154 & n1248;
  assign n5298 = ~n667 & n5297;
  assign n5299 = ~n278 & n5298;
  assign n5300 = ~n589 & n5299;
  assign n5301 = ~n712 & n5300;
  assign n5302 = ~n338 & n5301;
  assign n5303 = ~n564 & n5302;
  assign n5304 = ~n358 & n5303;
  assign n5305 = n2627 & n3264;
  assign n5306 = n3312 & n5305;
  assign n5307 = n5304 & n5306;
  assign n5308 = n1577 & n5307;
  assign n5309 = n247 & n5308;
  assign n5310 = n5296 & n5309;
  assign n5311 = n1254 & n5310;
  assign n5312 = n615 & n5311;
  assign n5313 = n5286 & n5312;
  assign n5314 = n100 & n5313;
  assign n5315 = ~n335 & n5314;
  assign n5316 = ~n402 & n5315;
  assign n5317 = ~n825 & n5316;
  assign n5318 = ~n296 & n5317;
  assign n5319 = ~n192 & n5318;
  assign n5320 = ~n429 & n5319;
  assign n5321 = ~n5254 & ~n5320;
  assign n5322 = n5254 & n5320;
  assign n5323 = ~n5321 & ~n5322;
  assign n5324 = ~ a[8]  & n5323;
  assign n5325 = ~n5321 & ~n5324;
  assign n5326 = n5053 & ~n5325;
  assign n5327 = n2880 & ~n2882;
  assign n5328 = ~n2883 & ~n5327;
  assign n5329 = n75 & n5328;
  assign n5330 = ~n1665 & n3020;
  assign n5331 = ~n1877 & n3023;
  assign n5332 = ~n1779 & n3028;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = ~n5330 & n5333;
  assign n5335 = ~n5329 & n5334;
  assign n5336 = ~n5053 & n5325;
  assign n5337 = ~n5326 & ~n5336;
  assign n5338 = ~n5335 & n5337;
  assign n5339 = ~n5326 & ~n5338;
  assign n5340 = ~n5169 & ~n5339;
  assign n5341 = ~n5170 & n5340;
  assign n5342 = ~n5169 & ~n5341;
  assign n5343 = n5134 & n5143;
  assign n5344 = ~n5144 & ~n5343;
  assign n5345 = ~n5342 & n5344;
  assign n5346 = ~n5144 & ~n5345;
  assign n5347 = ~n5131 & ~n5346;
  assign n5348 = n5131 & n5346;
  assign n5349 = ~n5347 & ~n5348;
  assign n5350 = ~n1060 & n3457;
  assign n5351 = ~n1235 & n3542;
  assign n5352 = ~n1178 & n3606;
  assign n5353 = ~n5351 & ~n5352;
  assign n5354 = ~n5350 & n5353;
  assign n5355 = ~n3368 & n5354;
  assign n5356 = ~n4429 & n5354;
  assign n5357 = ~n5355 & ~n5356;
  assign n5358 =  a[29]  & ~n5357;
  assign n5359 = ~ a[29]  & n5357;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = n5349 & ~n5360;
  assign n5362 = ~n5347 & ~n5361;
  assign n5363 = n5128 & ~n5362;
  assign n5364 = ~n5126 & ~n5363;
  assign n5365 = ~n4998 & ~n5364;
  assign n5366 = ~n4995 & ~n5365;
  assign n5367 = ~n4875 & n4886;
  assign n5368 = ~n4887 & ~n5367;
  assign n5369 = ~n5366 & n5368;
  assign n5370 = n5366 & ~n5368;
  assign n5371 = ~n5369 & ~n5370;
  assign n5372 = ~n3012 & n3884;
  assign n5373 = ~n587 & n3967;
  assign n5374 = ~n392 & n4046;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = ~n5372 & n5375;
  assign n5377 = n3018 & n4050;
  assign n5378 = n5376 & ~n5377;
  assign n5379 =  a[26]  & ~n5378;
  assign n5380 =  a[26]  & ~n5379;
  assign n5381 = ~n5378 & ~n5379;
  assign n5382 = ~n5380 & ~n5381;
  assign n5383 = n5371 & ~n5382;
  assign n5384 = ~n5369 & ~n5383;
  assign n5385 = ~n4980 & ~n5384;
  assign n5386 = n4980 & n5384;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = ~n3805 & n4694;
  assign n5389 = ~n3605 & n4533;
  assign n5390 = ~n3456 & n4604;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = ~n5388 & n5391;
  assign n5393 = n3818 & n4536;
  assign n5394 = n5392 & ~n5393;
  assign n5395 =  a[23]  & ~n5394;
  assign n5396 =  a[23]  & ~n5395;
  assign n5397 = ~n5394 & ~n5395;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = n5387 & ~n5398;
  assign n5400 = ~n5385 & ~n5399;
  assign n5401 = ~n4977 & ~n5400;
  assign n5402 = ~n4974 & ~n5401;
  assign n5403 = ~n4960 & ~n5402;
  assign n5404 = n4960 & n5402;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~n3877 & n4935;
  assign n5407 = ~n4927 & n4933;
  assign n5408 = ~n4515 & n5407;
  assign n5409 = ~n5406 & ~n5408;
  assign n5410 = n4609 & n4938;
  assign n5411 = n5409 & ~n5410;
  assign n5412 =  a[20]  & ~n5411;
  assign n5413 =  a[20]  & ~n5412;
  assign n5414 = ~n5411 & ~n5412;
  assign n5415 = ~n5413 & ~n5414;
  assign n5416 = n5405 & ~n5415;
  assign n5417 = ~n5403 & ~n5416;
  assign n5418 = ~n4957 & ~n5417;
  assign n5419 = n4957 & n5417;
  assign n5420 = ~n5418 & ~n5419;
  assign n5421 = n5405 & ~n5416;
  assign n5422 = ~n5415 & ~n5416;
  assign n5423 = ~n5421 & ~n5422;
  assign n5424 = n5387 & ~n5399;
  assign n5425 = ~n5398 & ~n5399;
  assign n5426 = ~n5424 & ~n5425;
  assign n5427 = n5371 & ~n5383;
  assign n5428 = ~n5382 & ~n5383;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = n4998 & n5364;
  assign n5431 = ~n5365 & ~n5430;
  assign n5432 = ~n392 & n3884;
  assign n5433 = ~n710 & n3967;
  assign n5434 = ~n587 & n4046;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = ~n5432 & n5435;
  assign n5437 = ~n4050 & n5436;
  assign n5438 = ~n3347 & n5436;
  assign n5439 = ~n5437 & ~n5438;
  assign n5440 =  a[26]  & ~n5439;
  assign n5441 = ~ a[26]  & n5439;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = n5431 & ~n5442;
  assign n5444 = ~n587 & n3884;
  assign n5445 = ~n867 & n3967;
  assign n5446 = ~n710 & n4046;
  assign n5447 = ~n5445 & ~n5446;
  assign n5448 = ~n5444 & n5447;
  assign n5449 = n3331 & n4050;
  assign n5450 = n5448 & ~n5449;
  assign n5451 =  a[26]  & ~n5450;
  assign n5452 =  a[26]  & ~n5451;
  assign n5453 = ~n5450 & ~n5451;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = ~n5128 & n5362;
  assign n5456 = ~n5363 & ~n5455;
  assign n5457 = ~n958 & n3457;
  assign n5458 = ~n1178 & n3542;
  assign n5459 = ~n1060 & n3606;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = ~n5457 & n5460;
  assign n5462 = ~n3368 & n5461;
  assign n5463 = ~n4633 & n5461;
  assign n5464 = ~n5462 & ~n5463;
  assign n5465 =  a[29]  & ~n5464;
  assign n5466 = ~ a[29]  & n5464;
  assign n5467 = ~n5465 & ~n5466;
  assign n5468 = n5456 & ~n5467;
  assign n5469 = ~n5456 & n5467;
  assign n5470 = ~n5468 & ~n5469;
  assign n5471 = ~n5454 & n5470;
  assign n5472 = ~n5468 & ~n5471;
  assign n5473 = ~n5431 & n5442;
  assign n5474 = ~n5443 & ~n5473;
  assign n5475 = ~n5472 & n5474;
  assign n5476 = ~n5443 & ~n5475;
  assign n5477 = ~n5429 & ~n5476;
  assign n5478 = n5429 & n5476;
  assign n5479 = ~n5477 & ~n5478;
  assign n5480 = ~n3456 & n4694;
  assign n5481 = ~n3539 & n4533;
  assign n5482 = ~n3605 & n4604;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = ~n5480 & n5483;
  assign n5485 = n3627 & n4536;
  assign n5486 = n5484 & ~n5485;
  assign n5487 =  a[23]  & ~n5486;
  assign n5488 =  a[23]  & ~n5487;
  assign n5489 = ~n5486 & ~n5487;
  assign n5490 = ~n5488 & ~n5489;
  assign n5491 = n5479 & ~n5490;
  assign n5492 = ~n5477 & ~n5491;
  assign n5493 = ~n5426 & ~n5492;
  assign n5494 = n5426 & n5492;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = n4930 & ~n4933;
  assign n5497 = ~n3877 & n5496;
  assign n5498 = ~n3964 & n4935;
  assign n5499 = ~n4045 & n5407;
  assign n5500 = ~n5498 & ~n5499;
  assign n5501 = ~n5497 & n5500;
  assign n5502 = n4067 & n4938;
  assign n5503 = n5501 & ~n5502;
  assign n5504 =  a[20]  & ~n5503;
  assign n5505 =  a[20]  & ~n5504;
  assign n5506 = ~n5503 & ~n5504;
  assign n5507 = ~n5505 & ~n5506;
  assign n5508 = n5495 & ~n5507;
  assign n5509 = ~n5493 & ~n5508;
  assign n5510 = ~n4515 & n5496;
  assign n5511 = ~n4045 & n4935;
  assign n5512 = ~n3877 & n5407;
  assign n5513 = ~n5511 & ~n5512;
  assign n5514 = ~n5510 & n5513;
  assign n5515 = ~n4938 & n5514;
  assign n5516 = ~n4715 & n5514;
  assign n5517 = ~n5515 & ~n5516;
  assign n5518 =  a[20]  & ~n5517;
  assign n5519 = ~ a[20]  & n5517;
  assign n5520 = ~n5518 & ~n5519;
  assign n5521 = ~n5509 & ~n5520;
  assign n5522 = n4977 & n5400;
  assign n5523 = ~n5401 & ~n5522;
  assign n5524 = n5509 & n5520;
  assign n5525 = ~n5521 & ~n5524;
  assign n5526 = n5523 & n5525;
  assign n5527 = ~n5521 & ~n5526;
  assign n5528 = ~n5423 & ~n5527;
  assign n5529 = n5423 & n5527;
  assign n5530 = ~n5528 & ~n5529;
  assign n5531 = n5479 & ~n5491;
  assign n5532 = ~n5490 & ~n5491;
  assign n5533 = ~n5531 & ~n5532;
  assign n5534 = ~n3605 & n4694;
  assign n5535 = ~n3012 & n4533;
  assign n5536 = ~n3539 & n4604;
  assign n5537 = ~n5535 & ~n5536;
  assign n5538 = ~n5534 & n5537;
  assign n5539 = n4084 & n4536;
  assign n5540 = n5538 & ~n5539;
  assign n5541 =  a[23]  & ~n5540;
  assign n5542 = ~n5540 & ~n5541;
  assign n5543 =  a[23]  & ~n5541;
  assign n5544 = ~n5542 & ~n5543;
  assign n5545 = n5472 & ~n5474;
  assign n5546 = ~n5475 & ~n5545;
  assign n5547 = ~n5544 & n5546;
  assign n5548 = ~n5544 & ~n5547;
  assign n5549 = n5546 & ~n5547;
  assign n5550 = ~n5548 & ~n5549;
  assign n5551 = n5470 & ~n5471;
  assign n5552 = ~n5454 & ~n5471;
  assign n5553 = ~n5551 & ~n5552;
  assign n5554 = ~n5339 & ~n5341;
  assign n5555 = ~n5170 & n5342;
  assign n5556 = ~n5554 & ~n5555;
  assign n5557 = ~n1572 & n3020;
  assign n5558 = ~n1665 & n3028;
  assign n5559 = ~n1779 & n3023;
  assign n5560 = n2884 & ~n2886;
  assign n5561 = ~n2887 & ~n5560;
  assign n5562 = n75 & n5561;
  assign n5563 = ~n5559 & ~n5562;
  assign n5564 = ~n5558 & n5563;
  assign n5565 = ~n5557 & n5564;
  assign n5566 = ~n5556 & ~n5565;
  assign n5567 = ~n1235 & n3457;
  assign n5568 = ~n1472 & n3542;
  assign n5569 = ~n1364 & n3606;
  assign n5570 = ~n5568 & ~n5569;
  assign n5571 = ~n5567 & n5570;
  assign n5572 = n3368 & n4848;
  assign n5573 = n5571 & ~n5572;
  assign n5574 =  a[29]  & ~n5573;
  assign n5575 = ~n5573 & ~n5574;
  assign n5576 =  a[29]  & ~n5574;
  assign n5577 = ~n5575 & ~n5576;
  assign n5578 = ~n5556 & ~n5566;
  assign n5579 = ~n5565 & ~n5566;
  assign n5580 = ~n5578 & ~n5579;
  assign n5581 = ~n5577 & ~n5580;
  assign n5582 = ~n5566 & ~n5581;
  assign n5583 = n5342 & ~n5344;
  assign n5584 = ~n5345 & ~n5583;
  assign n5585 = ~n5582 & n5584;
  assign n5586 = ~n1178 & n3457;
  assign n5587 = ~n1364 & n3542;
  assign n5588 = ~n1235 & n3606;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = ~n5586 & n5589;
  assign n5591 = n3368 & n4861;
  assign n5592 = n5590 & ~n5591;
  assign n5593 =  a[29]  & ~n5592;
  assign n5594 =  a[29]  & ~n5593;
  assign n5595 = ~n5592 & ~n5593;
  assign n5596 = ~n5594 & ~n5595;
  assign n5597 = n5582 & ~n5584;
  assign n5598 = ~n5585 & ~n5597;
  assign n5599 = ~n5596 & n5598;
  assign n5600 = ~n5585 & ~n5599;
  assign n5601 = ~n5349 & n5360;
  assign n5602 = ~n5361 & ~n5601;
  assign n5603 = ~n5600 & n5602;
  assign n5604 = n5600 & ~n5602;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = ~n710 & n3884;
  assign n5607 = ~n958 & n3967;
  assign n5608 = ~n867 & n4046;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = ~n5606 & n5609;
  assign n5611 = n4050 & n4179;
  assign n5612 = n5610 & ~n5611;
  assign n5613 =  a[26]  & ~n5612;
  assign n5614 =  a[26]  & ~n5613;
  assign n5615 = ~n5612 & ~n5613;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = n5605 & ~n5616;
  assign n5618 = ~n5603 & ~n5617;
  assign n5619 = ~n5553 & ~n5618;
  assign n5620 = n5553 & n5618;
  assign n5621 = ~n5619 & ~n5620;
  assign n5622 = ~n3539 & n4694;
  assign n5623 = ~n392 & n4533;
  assign n5624 = ~n3012 & n4604;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = ~n5622 & n5625;
  assign n5627 = n3715 & n4536;
  assign n5628 = n5626 & ~n5627;
  assign n5629 =  a[23]  & ~n5628;
  assign n5630 =  a[23]  & ~n5629;
  assign n5631 = ~n5628 & ~n5629;
  assign n5632 = ~n5630 & ~n5631;
  assign n5633 = n5621 & ~n5632;
  assign n5634 = ~n5619 & ~n5633;
  assign n5635 = ~n5550 & ~n5634;
  assign n5636 = ~n5547 & ~n5635;
  assign n5637 = ~n5533 & ~n5636;
  assign n5638 = n5533 & n5636;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = ~n4045 & n5496;
  assign n5641 = ~n3805 & n4935;
  assign n5642 = ~n3964 & n5407;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = ~n5640 & n5643;
  assign n5645 = n4477 & n4938;
  assign n5646 = n5644 & ~n5645;
  assign n5647 =  a[20]  & ~n5646;
  assign n5648 =  a[20]  & ~n5647;
  assign n5649 = ~n5646 & ~n5647;
  assign n5650 = ~n5648 & ~n5649;
  assign n5651 = n5639 & ~n5650;
  assign n5652 = ~n5637 & ~n5651;
  assign n5653 = ~ a[15]  &  a[16] ;
  assign n5654 =  a[15]  & ~ a[16] ;
  assign n5655 = ~n5653 & ~n5654;
  assign n5656 =  a[14]  & ~ a[15] ;
  assign n5657 = ~ a[14]  &  a[15] ;
  assign n5658 = ~n5656 & ~n5657;
  assign n5659 =  a[16]  & ~ a[17] ;
  assign n5660 = ~ a[16]  &  a[17] ;
  assign n5661 = ~n5659 & ~n5660;
  assign n5662 = n5658 & ~n5661;
  assign n5663 = n5655 & n5662;
  assign n5664 = ~n4515 & n5663;
  assign n5665 = ~n4522 & ~n5664;
  assign n5666 = ~n5658 & ~n5661;
  assign n5667 = ~n5664 & ~n5666;
  assign n5668 = ~n5665 & ~n5667;
  assign n5669 =  a[17]  & ~n5668;
  assign n5670 = ~ a[17]  & n5668;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = ~n5652 & ~n5671;
  assign n5673 = n5495 & ~n5508;
  assign n5674 = ~n5507 & ~n5508;
  assign n5675 = ~n5673 & ~n5674;
  assign n5676 = n5652 & n5671;
  assign n5677 = ~n5672 & ~n5676;
  assign n5678 = ~n5675 & n5677;
  assign n5679 = ~n5672 & ~n5678;
  assign n5680 = ~n5523 & ~n5525;
  assign n5681 = ~n5526 & ~n5680;
  assign n5682 = ~n5679 & n5681;
  assign n5683 = ~n5675 & ~n5678;
  assign n5684 = n5677 & ~n5678;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = n5639 & ~n5651;
  assign n5687 = ~n5650 & ~n5651;
  assign n5688 = ~n5686 & ~n5687;
  assign n5689 = n5550 & n5634;
  assign n5690 = ~n5635 & ~n5689;
  assign n5691 = ~n3964 & n5496;
  assign n5692 = ~n3456 & n4935;
  assign n5693 = ~n3805 & n5407;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = ~n5691 & n5694;
  assign n5696 = ~n4938 & n5695;
  assign n5697 = ~n4558 & n5695;
  assign n5698 = ~n5696 & ~n5697;
  assign n5699 =  a[20]  & ~n5698;
  assign n5700 = ~ a[20]  & n5698;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = n5690 & ~n5701;
  assign n5703 = n5621 & ~n5633;
  assign n5704 = ~n5632 & ~n5633;
  assign n5705 = ~n5703 & ~n5704;
  assign n5706 = n5605 & ~n5617;
  assign n5707 = ~n5616 & ~n5617;
  assign n5708 = ~n5706 & ~n5707;
  assign n5709 = n5598 & ~n5599;
  assign n5710 = ~n5596 & ~n5599;
  assign n5711 = ~n5709 & ~n5710;
  assign n5712 = ~n867 & n3884;
  assign n5713 = ~n1060 & n3967;
  assign n5714 = ~n958 & n4046;
  assign n5715 = ~n5713 & ~n5714;
  assign n5716 = ~n5712 & n5715;
  assign n5717 = ~n4050 & n5716;
  assign n5718 = ~n4204 & n5716;
  assign n5719 = ~n5717 & ~n5718;
  assign n5720 =  a[26]  & ~n5719;
  assign n5721 = ~ a[26]  & n5719;
  assign n5722 = ~n5720 & ~n5721;
  assign n5723 = ~n5711 & ~n5722;
  assign n5724 = ~n5577 & ~n5581;
  assign n5725 = ~n5580 & ~n5581;
  assign n5726 = ~n5724 & ~n5725;
  assign n5727 = ~n5335 & ~n5338;
  assign n5728 = n5337 & ~n5338;
  assign n5729 = ~n5727 & ~n5728;
  assign n5730 = ~ a[8]  & ~n5324;
  assign n5731 = ~n5322 & n5325;
  assign n5732 = ~n5730 & ~n5731;
  assign n5733 = n533 & n591;
  assign n5734 = ~n296 & n5733;
  assign n5735 = n3687 & n5734;
  assign n5736 = n3583 & n5735;
  assign n5737 = n1424 & n5736;
  assign n5738 = n3160 & n5737;
  assign n5739 = n977 & n5738;
  assign n5740 = n1575 & n5739;
  assign n5741 = ~n469 & n5740;
  assign n5742 = ~n884 & n5741;
  assign n5743 = ~n537 & n5742;
  assign n5744 = ~n1203 & n5743;
  assign n5745 = ~n449 & n5744;
  assign n5746 = ~n655 & n5745;
  assign n5747 = ~n289 & ~n364;
  assign n5748 = ~n287 & n5747;
  assign n5749 = n658 & n5748;
  assign n5750 = n5269 & n5749;
  assign n5751 = n824 & n5750;
  assign n5752 = n5239 & n5751;
  assign n5753 = n3205 & n5752;
  assign n5754 = n5746 & n5753;
  assign n5755 = n2633 & n5754;
  assign n5756 = n108 & n5755;
  assign n5757 = n570 & n5756;
  assign n5758 = ~n354 & n5757;
  assign n5759 = ~n115 & n5758;
  assign n5760 = ~n177 & n5759;
  assign n5761 = ~n357 & n5760;
  assign n5762 = ~n563 & n5761;
  assign n5763 = ~n173 & n5762;
  assign n5764 = ~n601 & n5763;
  assign n5765 = ~n283 & n5764;
  assign n5766 = n5254 & ~n5765;
  assign n5767 = ~n5254 & n5765;
  assign n5768 = n1497 & n3524;
  assign n5769 = ~n236 & n5768;
  assign n5770 = ~n504 & n5769;
  assign n5771 = ~n205 & n5770;
  assign n5772 = ~n537 & n5771;
  assign n5773 = ~n666 & n5772;
  assign n5774 = ~n364 & ~n430;
  assign n5775 = ~n127 & n5774;
  assign n5776 = ~n281 & ~n328;
  assign n5777 = ~n203 & n5776;
  assign n5778 = n5775 & n5777;
  assign n5779 = ~n242 & n5778;
  assign n5780 = ~n168 & n5779;
  assign n5781 = ~n884 & n5780;
  assign n5782 = ~n287 & n5781;
  assign n5783 = ~n961 & n5782;
  assign n5784 = ~n86 & n5783;
  assign n5785 = ~n158 & n5784;
  assign n5786 = ~n451 & ~n932;
  assign n5787 = ~n363 & n5786;
  assign n5788 = ~n136 & n5787;
  assign n5789 = ~n511 & n5788;
  assign n5790 = ~n275 & n5789;
  assign n5791 = ~n228 & n5790;
  assign n5792 = ~n151 & ~n602;
  assign n5793 = ~n189 & n5792;
  assign n5794 = n5791 & n5793;
  assign n5795 = n5785 & n5794;
  assign n5796 = n1237 & n5795;
  assign n5797 = n227 & n5796;
  assign n5798 = n100 & n5797;
  assign n5799 = n2758 & n5798;
  assign n5800 = ~n620 & n5799;
  assign n5801 = ~n506 & n5800;
  assign n5802 = ~n121 & n5801;
  assign n5803 = ~n527 & n5802;
  assign n5804 = ~n144 & n5803;
  assign n5805 = ~n493 & n5804;
  assign n5806 = ~n1127 & n5805;
  assign n5807 = ~n330 & ~n449;
  assign n5808 = ~n222 & n5807;
  assign n5809 = n2990 & n5808;
  assign n5810 = n5806 & n5809;
  assign n5811 = n4388 & n5810;
  assign n5812 = n616 & n5811;
  assign n5813 = n5773 & n5812;
  assign n5814 = n2651 & n5813;
  assign n5815 = n2940 & n5814;
  assign n5816 = n520 & n5815;
  assign n5817 = ~n847 & n5816;
  assign n5818 = ~n713 & n5817;
  assign n5819 = ~n171 & n5818;
  assign n5820 = ~n460 & n5819;
  assign n5821 = ~n331 & n5820;
  assign n5822 = ~n246 & n5821;
  assign n5823 = ~n623 & n5822;
  assign n5824 = ~n81 & n5823;
  assign n5825 = ~n231 & n5824;
  assign n5826 = ~ a[2]  & ~n5825;
  assign n5827 =  a[2]  & ~n5825;
  assign n5828 = ~ a[2]  & n5825;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = ~ a[5]  & ~n5829;
  assign n5831 = ~n5826 & ~n5830;
  assign n5832 = n5254 & ~n5831;
  assign n5833 = n2868 & ~n2870;
  assign n5834 = ~n2871 & ~n5833;
  assign n5835 = n75 & n5834;
  assign n5836 = ~n1913 & n3020;
  assign n5837 = ~n2057 & n3023;
  assign n5838 = ~n1992 & n3028;
  assign n5839 = ~n5837 & ~n5838;
  assign n5840 = ~n5836 & n5839;
  assign n5841 = ~n5835 & n5840;
  assign n5842 = ~n5254 & n5831;
  assign n5843 = ~n5832 & ~n5842;
  assign n5844 = ~n5841 & n5843;
  assign n5845 = ~n5832 & ~n5844;
  assign n5846 = ~n5766 & ~n5845;
  assign n5847 = ~n5767 & n5846;
  assign n5848 = ~n5766 & ~n5847;
  assign n5849 = ~n5732 & ~n5848;
  assign n5850 = n2876 & ~n2878;
  assign n5851 = ~n2879 & ~n5850;
  assign n5852 = n75 & n5851;
  assign n5853 = ~n1779 & n3020;
  assign n5854 = ~n1913 & n3023;
  assign n5855 = ~n1877 & n3028;
  assign n5856 = ~n5854 & ~n5855;
  assign n5857 = ~n5853 & n5856;
  assign n5858 = ~n5852 & n5857;
  assign n5859 = n5732 & n5848;
  assign n5860 = ~n5849 & ~n5859;
  assign n5861 = ~n5858 & n5860;
  assign n5862 = ~n5849 & ~n5861;
  assign n5863 = ~n5729 & ~n5862;
  assign n5864 = n5729 & n5862;
  assign n5865 = ~n5863 & ~n5864;
  assign n5866 = ~n1364 & n3457;
  assign n5867 = ~n1572 & n3542;
  assign n5868 = ~n1472 & n3606;
  assign n5869 = ~n5867 & ~n5868;
  assign n5870 = ~n5866 & n5869;
  assign n5871 = ~n3368 & n5870;
  assign n5872 = ~n5114 & n5870;
  assign n5873 = ~n5871 & ~n5872;
  assign n5874 =  a[29]  & ~n5873;
  assign n5875 = ~ a[29]  & n5873;
  assign n5876 = ~n5874 & ~n5875;
  assign n5877 = n5865 & ~n5876;
  assign n5878 = ~n5863 & ~n5877;
  assign n5879 = ~n5726 & ~n5878;
  assign n5880 = n5726 & n5878;
  assign n5881 = ~n5879 & ~n5880;
  assign n5882 = ~n958 & n3884;
  assign n5883 = ~n1178 & n3967;
  assign n5884 = ~n1060 & n4046;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = ~n5882 & n5885;
  assign n5887 = n4050 & n4633;
  assign n5888 = n5886 & ~n5887;
  assign n5889 =  a[26]  & ~n5888;
  assign n5890 =  a[26]  & ~n5889;
  assign n5891 = ~n5888 & ~n5889;
  assign n5892 = ~n5890 & ~n5891;
  assign n5893 = n5881 & ~n5892;
  assign n5894 = ~n5879 & ~n5893;
  assign n5895 = n5711 & n5722;
  assign n5896 = ~n5723 & ~n5895;
  assign n5897 = ~n5894 & n5896;
  assign n5898 = ~n5723 & ~n5897;
  assign n5899 = ~n5708 & ~n5898;
  assign n5900 = n5708 & n5898;
  assign n5901 = ~n5899 & ~n5900;
  assign n5902 = ~n3012 & n4694;
  assign n5903 = ~n587 & n4533;
  assign n5904 = ~n392 & n4604;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = ~n5902 & n5905;
  assign n5907 = n3018 & n4536;
  assign n5908 = n5906 & ~n5907;
  assign n5909 =  a[23]  & ~n5908;
  assign n5910 =  a[23]  & ~n5909;
  assign n5911 = ~n5908 & ~n5909;
  assign n5912 = ~n5910 & ~n5911;
  assign n5913 = n5901 & ~n5912;
  assign n5914 = ~n5899 & ~n5913;
  assign n5915 = ~n5705 & ~n5914;
  assign n5916 = n5705 & n5914;
  assign n5917 = ~n5915 & ~n5916;
  assign n5918 = ~n3805 & n5496;
  assign n5919 = ~n3605 & n4935;
  assign n5920 = ~n3456 & n5407;
  assign n5921 = ~n5919 & ~n5920;
  assign n5922 = ~n5918 & n5921;
  assign n5923 = n3818 & n4938;
  assign n5924 = n5922 & ~n5923;
  assign n5925 =  a[20]  & ~n5924;
  assign n5926 =  a[20]  & ~n5925;
  assign n5927 = ~n5924 & ~n5925;
  assign n5928 = ~n5926 & ~n5927;
  assign n5929 = n5917 & ~n5928;
  assign n5930 = ~n5915 & ~n5929;
  assign n5931 = ~n5690 & n5701;
  assign n5932 = ~n5702 & ~n5931;
  assign n5933 = ~n5930 & n5932;
  assign n5934 = ~n5702 & ~n5933;
  assign n5935 = ~n5688 & ~n5934;
  assign n5936 = n5688 & n5934;
  assign n5937 = ~n5935 & ~n5936;
  assign n5938 = ~n3877 & n5663;
  assign n5939 = ~n5655 & n5658;
  assign n5940 = ~n4515 & n5939;
  assign n5941 = ~n5938 & ~n5940;
  assign n5942 = n4609 & n5666;
  assign n5943 = n5941 & ~n5942;
  assign n5944 =  a[17]  & ~n5943;
  assign n5945 =  a[17]  & ~n5944;
  assign n5946 = ~n5943 & ~n5944;
  assign n5947 = ~n5945 & ~n5946;
  assign n5948 = n5937 & ~n5947;
  assign n5949 = ~n5935 & ~n5948;
  assign n5950 = ~n5685 & ~n5949;
  assign n5951 = n5685 & n5949;
  assign n5952 = ~n5950 & ~n5951;
  assign n5953 = n5937 & ~n5948;
  assign n5954 = ~n5947 & ~n5948;
  assign n5955 = ~n5953 & ~n5954;
  assign n5956 = n5917 & ~n5929;
  assign n5957 = ~n5928 & ~n5929;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = n5901 & ~n5913;
  assign n5960 = ~n5912 & ~n5913;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = ~n392 & n4694;
  assign n5963 = ~n710 & n4533;
  assign n5964 = ~n587 & n4604;
  assign n5965 = ~n5963 & ~n5964;
  assign n5966 = ~n5962 & n5965;
  assign n5967 = n3347 & n4536;
  assign n5968 = n5966 & ~n5967;
  assign n5969 =  a[23]  & ~n5968;
  assign n5970 = ~n5968 & ~n5969;
  assign n5971 =  a[23]  & ~n5969;
  assign n5972 = ~n5970 & ~n5971;
  assign n5973 = n5894 & ~n5896;
  assign n5974 = ~n5897 & ~n5973;
  assign n5975 = ~n5972 & n5974;
  assign n5976 = ~n5972 & ~n5975;
  assign n5977 = n5974 & ~n5975;
  assign n5978 = ~n5976 & ~n5977;
  assign n5979 = n5881 & ~n5893;
  assign n5980 = ~n5892 & ~n5893;
  assign n5981 = ~n5979 & ~n5980;
  assign n5982 = ~n1472 & n3457;
  assign n5983 = ~n1665 & n3542;
  assign n5984 = ~n1572 & n3606;
  assign n5985 = ~n5983 & ~n5984;
  assign n5986 = ~n5982 & n5985;
  assign n5987 = n3368 & n5139;
  assign n5988 = n5986 & ~n5987;
  assign n5989 =  a[29]  & ~n5988;
  assign n5990 = ~n5988 & ~n5989;
  assign n5991 =  a[29]  & ~n5989;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = ~n5858 & ~n5861;
  assign n5994 = n5860 & ~n5861;
  assign n5995 = ~n5993 & ~n5994;
  assign n5996 = ~n5992 & ~n5995;
  assign n5997 = ~n5992 & ~n5996;
  assign n5998 = ~n5995 & ~n5996;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = ~n5845 & ~n5847;
  assign n6001 = ~n5767 & n5848;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~n1877 & n3020;
  assign n6004 = ~n1913 & n3028;
  assign n6005 = ~n1992 & n3023;
  assign n6006 = n2872 & ~n2874;
  assign n6007 = ~n2875 & ~n6006;
  assign n6008 = n75 & n6007;
  assign n6009 = ~n6005 & ~n6008;
  assign n6010 = ~n6004 & n6009;
  assign n6011 = ~n6003 & n6010;
  assign n6012 = ~n6002 & ~n6011;
  assign n6013 = ~n5841 & ~n5844;
  assign n6014 = n5843 & ~n5844;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = ~n289 & n2059;
  assign n6017 = ~n620 & n6016;
  assign n6018 = ~n352 & n6017;
  assign n6019 = ~n394 & n6018;
  assign n6020 = ~n603 & n6019;
  assign n6021 = n1727 & n2705;
  assign n6022 = n2556 & n6021;
  assign n6023 = ~n330 & n6022;
  assign n6024 = ~n466 & n6023;
  assign n6025 = n1680 & n6024;
  assign n6026 = ~n270 & n6025;
  assign n6027 = n4335 & n5152;
  assign n6028 = n5056 & n6027;
  assign n6029 = n1084 & n6028;
  assign n6030 = n2127 & n6029;
  assign n6031 = n3580 & n6030;
  assign n6032 = n6026 & n6031;
  assign n6033 = n2439 & n6032;
  assign n6034 = n6020 & n6033;
  assign n6035 = n1029 & n6034;
  assign n6036 = n4786 & n6035;
  assign n6037 = n618 & n6036;
  assign n6038 = ~n243 & n6037;
  assign n6039 = ~n519 & n6038;
  assign n6040 = ~n127 & n6039;
  assign n6041 = ~n81 & n6040;
  assign n6042 =  a[2]  & ~n6041;
  assign n6043 = ~ a[2]  & n6041;
  assign n6044 = n467 & n1611;
  assign n6045 = ~n420 & n6044;
  assign n6046 = ~n1062 & n6045;
  assign n6047 = ~n417 & n6046;
  assign n6048 = ~n400 & n6047;
  assign n6049 = ~n416 & n6048;
  assign n6050 = ~n192 & n6049;
  assign n6051 = ~n563 & n6050;
  assign n6052 = ~n425 & n6051;
  assign n6053 = ~n714 & n6052;
  assign n6054 = ~n243 & n6053;
  assign n6055 = n690 & n3252;
  assign n6056 = n618 & n6055;
  assign n6057 = n4828 & n6056;
  assign n6058 = n204 & n6057;
  assign n6059 = n324 & n6058;
  assign n6060 = n6054 & n6059;
  assign n6061 = n2623 & n6060;
  assign n6062 = n2961 & n6061;
  assign n6063 = n4274 & n6062;
  assign n6064 = n604 & n6063;
  assign n6065 = n454 & n6064;
  assign n6066 = n423 & n6065;
  assign n6067 = n731 & n6066;
  assign n6068 = n1379 & n6067;
  assign n6069 = ~n149 & n6068;
  assign n6070 = ~n246 & n6069;
  assign n6071 = ~n791 & n6070;
  assign n6072 = ~n592 & n6071;
  assign n6073 = ~n886 & n6072;
  assign n6074 = ~n449 & n6073;
  assign n6075 =  a[2]  & ~n6074;
  assign n6076 = ~ a[2]  & n6074;
  assign n6077 = n1426 & n1644;
  assign n6078 = ~n190 & n6077;
  assign n6079 = ~n239 & n6078;
  assign n6080 = ~n637 & n6079;
  assign n6081 = ~n305 & n6080;
  assign n6082 = ~n130 & n6081;
  assign n6083 = ~n1010 & n6082;
  assign n6084 = ~n295 & ~n395;
  assign n6085 = n2593 & n5150;
  assign n6086 = n1438 & n6085;
  assign n6087 = n6084 & n6086;
  assign n6088 = n5193 & n6087;
  assign n6089 = n1601 & n6088;
  assign n6090 = n1029 & n6089;
  assign n6091 = n454 & n6090;
  assign n6092 = n979 & n6091;
  assign n6093 = ~n752 & n6092;
  assign n6094 = ~n224 & n6093;
  assign n6095 = ~n275 & n6094;
  assign n6096 = ~n226 & n6095;
  assign n6097 = ~n451 & n6096;
  assign n6098 = n590 & ~n1072;
  assign n6099 = ~n206 & n6098;
  assign n6100 = ~n714 & n6099;
  assign n6101 = ~n689 & n6100;
  assign n6102 = ~n474 & n6101;
  assign n6103 = ~n111 & n4367;
  assign n6104 = ~n603 & n6103;
  assign n6105 = n4269 & n6104;
  assign n6106 = n2241 & n6105;
  assign n6107 = n2807 & n6106;
  assign n6108 = n6102 & n6107;
  assign n6109 = n2751 & n6108;
  assign n6110 = n6097 & n6109;
  assign n6111 = n6083 & n6110;
  assign n6112 = n333 & n6111;
  assign n6113 = n1291 & n6112;
  assign n6114 = n4786 & n6113;
  assign n6115 = ~n201 & n6114;
  assign n6116 = ~n564 & n6115;
  assign n6117 = ~n489 & n6116;
  assign n6118 = ~n886 & n6117;
  assign n6119 =  a[2]  & ~n6118;
  assign n6120 = ~ a[2]  & n6118;
  assign n6121 = n2852 & ~n2854;
  assign n6122 = ~n2855 & ~n6121;
  assign n6123 = n75 & n6122;
  assign n6124 = ~n2189 & n3020;
  assign n6125 = ~n2388 & n3023;
  assign n6126 = ~n2291 & n3028;
  assign n6127 = ~n6125 & ~n6126;
  assign n6128 = ~n6124 & n6127;
  assign n6129 = ~n6123 & n6128;
  assign n6130 = ~n6119 & ~n6129;
  assign n6131 = ~n6120 & n6130;
  assign n6132 = ~n6119 & ~n6131;
  assign n6133 = ~n6075 & ~n6132;
  assign n6134 = ~n6076 & n6133;
  assign n6135 = ~n6075 & ~n6134;
  assign n6136 = ~n6042 & ~n6135;
  assign n6137 = ~n6043 & n6136;
  assign n6138 = ~n6042 & ~n6137;
  assign n6139 =  a[5]  & n5829;
  assign n6140 = ~n5830 & ~n6139;
  assign n6141 = ~n6138 & n6140;
  assign n6142 = n2864 & ~n2866;
  assign n6143 = ~n2867 & ~n6142;
  assign n6144 = n75 & n6143;
  assign n6145 = ~n1992 & n3020;
  assign n6146 = ~n2152 & n3023;
  assign n6147 = ~n2057 & n3028;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = ~n6145 & n6148;
  assign n6150 = ~n6144 & n6149;
  assign n6151 = n6138 & ~n6140;
  assign n6152 = ~n6141 & ~n6151;
  assign n6153 = ~n6150 & n6152;
  assign n6154 = ~n6141 & ~n6153;
  assign n6155 = ~n6015 & ~n6154;
  assign n6156 = n6015 & n6154;
  assign n6157 = ~n6155 & ~n6156;
  assign n6158 = ~n1665 & n3457;
  assign n6159 = ~n1877 & n3542;
  assign n6160 = ~n1779 & n3606;
  assign n6161 = ~n6159 & ~n6160;
  assign n6162 = ~n6158 & n6161;
  assign n6163 = ~n3368 & n6162;
  assign n6164 = ~n5328 & n6162;
  assign n6165 = ~n6163 & ~n6164;
  assign n6166 =  a[29]  & ~n6165;
  assign n6167 = ~ a[29]  & n6165;
  assign n6168 = ~n6166 & ~n6167;
  assign n6169 = n6157 & ~n6168;
  assign n6170 = ~n6155 & ~n6169;
  assign n6171 = ~n6002 & ~n6012;
  assign n6172 = ~n6011 & ~n6012;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = ~n6170 & ~n6173;
  assign n6175 = ~n6012 & ~n6174;
  assign n6176 = ~n5999 & ~n6175;
  assign n6177 = ~n5996 & ~n6176;
  assign n6178 = ~n5865 & n5876;
  assign n6179 = ~n5877 & ~n6178;
  assign n6180 = ~n6177 & n6179;
  assign n6181 = n6177 & ~n6179;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = ~n1060 & n3884;
  assign n6184 = ~n1235 & n3967;
  assign n6185 = ~n1178 & n4046;
  assign n6186 = ~n6184 & ~n6185;
  assign n6187 = ~n6183 & n6186;
  assign n6188 = n4050 & n4429;
  assign n6189 = n6187 & ~n6188;
  assign n6190 =  a[26]  & ~n6189;
  assign n6191 =  a[26]  & ~n6190;
  assign n6192 = ~n6189 & ~n6190;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = n6182 & ~n6193;
  assign n6195 = ~n6180 & ~n6194;
  assign n6196 = ~n5981 & ~n6195;
  assign n6197 = n5981 & n6195;
  assign n6198 = ~n6196 & ~n6197;
  assign n6199 = ~n587 & n4694;
  assign n6200 = ~n867 & n4533;
  assign n6201 = ~n710 & n4604;
  assign n6202 = ~n6200 & ~n6201;
  assign n6203 = ~n6199 & n6202;
  assign n6204 = n3331 & n4536;
  assign n6205 = n6203 & ~n6204;
  assign n6206 =  a[23]  & ~n6205;
  assign n6207 =  a[23]  & ~n6206;
  assign n6208 = ~n6205 & ~n6206;
  assign n6209 = ~n6207 & ~n6208;
  assign n6210 = n6198 & ~n6209;
  assign n6211 = ~n6196 & ~n6210;
  assign n6212 = ~n5978 & ~n6211;
  assign n6213 = ~n5975 & ~n6212;
  assign n6214 = ~n5961 & ~n6213;
  assign n6215 = n5961 & n6213;
  assign n6216 = ~n6214 & ~n6215;
  assign n6217 = ~n3456 & n5496;
  assign n6218 = ~n3539 & n4935;
  assign n6219 = ~n3605 & n5407;
  assign n6220 = ~n6218 & ~n6219;
  assign n6221 = ~n6217 & n6220;
  assign n6222 = n3627 & n4938;
  assign n6223 = n6221 & ~n6222;
  assign n6224 =  a[20]  & ~n6223;
  assign n6225 =  a[20]  & ~n6224;
  assign n6226 = ~n6223 & ~n6224;
  assign n6227 = ~n6225 & ~n6226;
  assign n6228 = n6216 & ~n6227;
  assign n6229 = ~n6214 & ~n6228;
  assign n6230 = ~n5958 & ~n6229;
  assign n6231 = n5958 & n6229;
  assign n6232 = ~n6230 & ~n6231;
  assign n6233 = ~n5658 & n5661;
  assign n6234 = ~n3877 & n6233;
  assign n6235 = ~n3964 & n5663;
  assign n6236 = ~n4045 & n5939;
  assign n6237 = ~n6235 & ~n6236;
  assign n6238 = ~n6234 & n6237;
  assign n6239 = n4067 & n5666;
  assign n6240 = n6238 & ~n6239;
  assign n6241 =  a[17]  & ~n6240;
  assign n6242 =  a[17]  & ~n6241;
  assign n6243 = ~n6240 & ~n6241;
  assign n6244 = ~n6242 & ~n6243;
  assign n6245 = n6232 & ~n6244;
  assign n6246 = ~n6230 & ~n6245;
  assign n6247 = ~n4515 & n6233;
  assign n6248 = ~n4045 & n5663;
  assign n6249 = ~n3877 & n5939;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~n6247 & n6250;
  assign n6252 = ~n5666 & n6251;
  assign n6253 = ~n4715 & n6251;
  assign n6254 = ~n6252 & ~n6253;
  assign n6255 =  a[17]  & ~n6254;
  assign n6256 = ~ a[17]  & n6254;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = ~n6246 & ~n6257;
  assign n6259 = n6246 & n6257;
  assign n6260 = ~n6258 & ~n6259;
  assign n6261 = n5930 & ~n5932;
  assign n6262 = ~n5933 & ~n6261;
  assign n6263 = n6260 & n6262;
  assign n6264 = ~n6258 & ~n6263;
  assign n6265 = ~n5955 & ~n6264;
  assign n6266 = n5955 & n6264;
  assign n6267 = ~n6265 & ~n6266;
  assign n6268 = n6216 & ~n6228;
  assign n6269 = ~n6227 & ~n6228;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = n5978 & n6211;
  assign n6272 = ~n6212 & ~n6271;
  assign n6273 = ~n3605 & n5496;
  assign n6274 = ~n3012 & n4935;
  assign n6275 = ~n3539 & n5407;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = ~n6273 & n6276;
  assign n6278 = ~n4938 & n6277;
  assign n6279 = ~n4084 & n6277;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 =  a[20]  & ~n6280;
  assign n6282 = ~ a[20]  & n6280;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = n6272 & ~n6283;
  assign n6285 = n6198 & ~n6210;
  assign n6286 = ~n6209 & ~n6210;
  assign n6287 = ~n6285 & ~n6286;
  assign n6288 = n6182 & ~n6194;
  assign n6289 = ~n6193 & ~n6194;
  assign n6290 = ~n6288 & ~n6289;
  assign n6291 = n5999 & n6175;
  assign n6292 = ~n6176 & ~n6291;
  assign n6293 = ~n1178 & n3884;
  assign n6294 = ~n1364 & n3967;
  assign n6295 = ~n1235 & n4046;
  assign n6296 = ~n6294 & ~n6295;
  assign n6297 = ~n6293 & n6296;
  assign n6298 = ~n4050 & n6297;
  assign n6299 = ~n4861 & n6297;
  assign n6300 = ~n6298 & ~n6299;
  assign n6301 =  a[26]  & ~n6300;
  assign n6302 = ~ a[26]  & n6300;
  assign n6303 = ~n6301 & ~n6302;
  assign n6304 = n6292 & ~n6303;
  assign n6305 = ~n6170 & ~n6174;
  assign n6306 = ~n6173 & ~n6174;
  assign n6307 = ~n6305 & ~n6306;
  assign n6308 = ~n1572 & n3457;
  assign n6309 = ~n1779 & n3542;
  assign n6310 = ~n1665 & n3606;
  assign n6311 = ~n6309 & ~n6310;
  assign n6312 = ~n6308 & n6311;
  assign n6313 = ~n3368 & n6312;
  assign n6314 = ~n5561 & n6312;
  assign n6315 = ~n6313 & ~n6314;
  assign n6316 =  a[29]  & ~n6315;
  assign n6317 = ~ a[29]  & n6315;
  assign n6318 = ~n6316 & ~n6317;
  assign n6319 = ~n6307 & ~n6318;
  assign n6320 = n6307 & n6318;
  assign n6321 = ~n6319 & ~n6320;
  assign n6322 = ~n1235 & n3884;
  assign n6323 = ~n1472 & n3967;
  assign n6324 = ~n1364 & n4046;
  assign n6325 = ~n6323 & ~n6324;
  assign n6326 = ~n6322 & n6325;
  assign n6327 = n4050 & n4848;
  assign n6328 = n6326 & ~n6327;
  assign n6329 =  a[26]  & ~n6328;
  assign n6330 =  a[26]  & ~n6329;
  assign n6331 = ~n6328 & ~n6329;
  assign n6332 = ~n6330 & ~n6331;
  assign n6333 = n6321 & ~n6332;
  assign n6334 = ~n6319 & ~n6333;
  assign n6335 = ~n6292 & n6303;
  assign n6336 = ~n6304 & ~n6335;
  assign n6337 = ~n6334 & n6336;
  assign n6338 = ~n6304 & ~n6337;
  assign n6339 = ~n6290 & ~n6338;
  assign n6340 = n6290 & n6338;
  assign n6341 = ~n6339 & ~n6340;
  assign n6342 = ~n710 & n4694;
  assign n6343 = ~n958 & n4533;
  assign n6344 = ~n867 & n4604;
  assign n6345 = ~n6343 & ~n6344;
  assign n6346 = ~n6342 & n6345;
  assign n6347 = n4179 & n4536;
  assign n6348 = n6346 & ~n6347;
  assign n6349 =  a[23]  & ~n6348;
  assign n6350 =  a[23]  & ~n6349;
  assign n6351 = ~n6348 & ~n6349;
  assign n6352 = ~n6350 & ~n6351;
  assign n6353 = n6341 & ~n6352;
  assign n6354 = ~n6339 & ~n6353;
  assign n6355 = ~n6287 & ~n6354;
  assign n6356 = n6287 & n6354;
  assign n6357 = ~n6355 & ~n6356;
  assign n6358 = ~n3539 & n5496;
  assign n6359 = ~n392 & n4935;
  assign n6360 = ~n3012 & n5407;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = ~n6358 & n6361;
  assign n6363 = n3715 & n4938;
  assign n6364 = n6362 & ~n6363;
  assign n6365 =  a[20]  & ~n6364;
  assign n6366 =  a[20]  & ~n6365;
  assign n6367 = ~n6364 & ~n6365;
  assign n6368 = ~n6366 & ~n6367;
  assign n6369 = n6357 & ~n6368;
  assign n6370 = ~n6355 & ~n6369;
  assign n6371 = ~n6272 & n6283;
  assign n6372 = ~n6284 & ~n6371;
  assign n6373 = ~n6370 & n6372;
  assign n6374 = ~n6284 & ~n6373;
  assign n6375 = ~n6270 & ~n6374;
  assign n6376 = n6270 & n6374;
  assign n6377 = ~n6375 & ~n6376;
  assign n6378 = ~n4045 & n6233;
  assign n6379 = ~n3805 & n5663;
  assign n6380 = ~n3964 & n5939;
  assign n6381 = ~n6379 & ~n6380;
  assign n6382 = ~n6378 & n6381;
  assign n6383 = n4477 & n5666;
  assign n6384 = n6382 & ~n6383;
  assign n6385 =  a[17]  & ~n6384;
  assign n6386 =  a[17]  & ~n6385;
  assign n6387 = ~n6384 & ~n6385;
  assign n6388 = ~n6386 & ~n6387;
  assign n6389 = n6377 & ~n6388;
  assign n6390 = ~n6375 & ~n6389;
  assign n6391 =  a[11]  & ~ a[12] ;
  assign n6392 = ~ a[11]  &  a[12] ;
  assign n6393 = ~n6391 & ~n6392;
  assign n6394 =  a[13]  & ~ a[14] ;
  assign n6395 = ~ a[13]  &  a[14] ;
  assign n6396 = ~n6394 & ~n6395;
  assign n6397 = ~n6393 & ~n6396;
  assign n6398 = ~ a[12]  &  a[13] ;
  assign n6399 =  a[12]  & ~ a[13] ;
  assign n6400 = ~n6398 & ~n6399;
  assign n6401 = n6393 & ~n6396;
  assign n6402 = n6400 & n6401;
  assign n6403 = ~n4515 & n6402;
  assign n6404 = ~n6397 & ~n6403;
  assign n6405 = ~n4522 & ~n6403;
  assign n6406 = ~n6404 & ~n6405;
  assign n6407 =  a[14]  & ~n6406;
  assign n6408 = ~ a[14]  & n6406;
  assign n6409 = ~n6407 & ~n6408;
  assign n6410 = ~n6390 & ~n6409;
  assign n6411 = n6232 & ~n6245;
  assign n6412 = ~n6244 & ~n6245;
  assign n6413 = ~n6411 & ~n6412;
  assign n6414 = n6390 & n6409;
  assign n6415 = ~n6410 & ~n6414;
  assign n6416 = ~n6413 & n6415;
  assign n6417 = ~n6410 & ~n6416;
  assign n6418 = ~n6260 & ~n6262;
  assign n6419 = ~n6263 & ~n6418;
  assign n6420 = ~n6417 & n6419;
  assign n6421 = n6417 & ~n6419;
  assign n6422 = ~n6420 & ~n6421;
  assign n6423 = ~n6413 & ~n6416;
  assign n6424 = n6415 & ~n6416;
  assign n6425 = ~n6423 & ~n6424;
  assign n6426 = ~n3964 & n6233;
  assign n6427 = ~n3456 & n5663;
  assign n6428 = ~n3805 & n5939;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = ~n6426 & n6429;
  assign n6431 = n4558 & n5666;
  assign n6432 = n6430 & ~n6431;
  assign n6433 =  a[17]  & ~n6432;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 =  a[17]  & ~n6433;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = n6370 & ~n6372;
  assign n6438 = ~n6373 & ~n6437;
  assign n6439 = ~n6436 & n6438;
  assign n6440 = ~n6436 & ~n6439;
  assign n6441 = n6438 & ~n6439;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = n6357 & ~n6369;
  assign n6444 = ~n6368 & ~n6369;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = n6341 & ~n6353;
  assign n6447 = ~n6352 & ~n6353;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = ~n867 & n4694;
  assign n6450 = ~n1060 & n4533;
  assign n6451 = ~n958 & n4604;
  assign n6452 = ~n6450 & ~n6451;
  assign n6453 = ~n6449 & n6452;
  assign n6454 = n4204 & n4536;
  assign n6455 = n6453 & ~n6454;
  assign n6456 =  a[23]  & ~n6455;
  assign n6457 = ~n6455 & ~n6456;
  assign n6458 =  a[23]  & ~n6456;
  assign n6459 = ~n6457 & ~n6458;
  assign n6460 = n6334 & ~n6336;
  assign n6461 = ~n6337 & ~n6460;
  assign n6462 = ~n6459 & n6461;
  assign n6463 = ~n6459 & ~n6462;
  assign n6464 = n6461 & ~n6462;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = n6321 & ~n6333;
  assign n6467 = ~n6332 & ~n6333;
  assign n6468 = ~n6466 & ~n6467;
  assign n6469 = n6152 & ~n6153;
  assign n6470 = ~n6150 & ~n6153;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = ~n6135 & ~n6137;
  assign n6473 = ~n6043 & n6138;
  assign n6474 = ~n6472 & ~n6473;
  assign n6475 = ~n2057 & n3020;
  assign n6476 = ~n2152 & n3028;
  assign n6477 = ~n2189 & n3023;
  assign n6478 = n2860 & ~n2862;
  assign n6479 = ~n2863 & ~n6478;
  assign n6480 = n75 & n6479;
  assign n6481 = ~n6477 & ~n6480;
  assign n6482 = ~n6476 & n6481;
  assign n6483 = ~n6475 & n6482;
  assign n6484 = ~n6474 & ~n6483;
  assign n6485 = ~n6132 & ~n6134;
  assign n6486 = ~n6076 & n6135;
  assign n6487 = ~n6485 & ~n6486;
  assign n6488 = ~n2152 & n3020;
  assign n6489 = ~n2189 & n3028;
  assign n6490 = ~n2291 & n3023;
  assign n6491 = n2856 & ~n2858;
  assign n6492 = ~n2859 & ~n6491;
  assign n6493 = n75 & n6492;
  assign n6494 = ~n6490 & ~n6493;
  assign n6495 = ~n6489 & n6494;
  assign n6496 = ~n6488 & n6495;
  assign n6497 = ~n6487 & ~n6496;
  assign n6498 = ~n6129 & ~n6131;
  assign n6499 = ~n6120 & n6132;
  assign n6500 = ~n6498 & ~n6499;
  assign n6501 = n2608 & n4357;
  assign n6502 = n4828 & n6501;
  assign n6503 = n4279 & n6502;
  assign n6504 = n1794 & n6503;
  assign n6505 = n1292 & n6504;
  assign n6506 = n874 & n6505;
  assign n6507 = n1139 & n6506;
  assign n6508 = n2993 & n6507;
  assign n6509 = n116 & n6508;
  assign n6510 = ~n617 & n6509;
  assign n6511 = ~n254 & n6510;
  assign n6512 = ~n809 & n6511;
  assign n6513 = ~n368 & n6512;
  assign n6514 = ~n791 & n6513;
  assign n6515 = ~n175 & n5171;
  assign n6516 = ~n206 & n6515;
  assign n6517 = ~n655 & n6516;
  assign n6518 = ~n123 & ~n518;
  assign n6519 = ~n157 & n6518;
  assign n6520 = ~n270 & n6519;
  assign n6521 = n3524 & n5775;
  assign n6522 = n691 & n6521;
  assign n6523 = n6520 & n6522;
  assign n6524 = n6517 & n6523;
  assign n6525 = n1709 & n6524;
  assign n6526 = n4405 & n6525;
  assign n6527 = n4375 & n6526;
  assign n6528 = n6514 & n6527;
  assign n6529 = n454 & n6528;
  assign n6530 = n731 & n6529;
  assign n6531 = n1478 & n6530;
  assign n6532 = ~n136 & n6531;
  assign n6533 = ~n248 & n6532;
  assign n6534 = ~n298 & n6533;
  assign n6535 = ~n273 & n6534;
  assign n6536 = ~n436 & n6535;
  assign n6537 = ~n2291 & n3020;
  assign n6538 = ~n2388 & n3028;
  assign n6539 = ~n2464 & n3023;
  assign n6540 = n2848 & ~n2850;
  assign n6541 = ~n2851 & ~n6540;
  assign n6542 = n75 & n6541;
  assign n6543 = ~n6539 & ~n6542;
  assign n6544 = ~n6538 & n6543;
  assign n6545 = ~n6537 & n6544;
  assign n6546 = ~n6536 & ~n6545;
  assign n6547 = ~n278 & ~n396;
  assign n6548 = ~n532 & n6547;
  assign n6549 = n5021 & n6548;
  assign n6550 = n1785 & n6549;
  assign n6551 = n1586 & n6550;
  assign n6552 = n4127 & n6551;
  assign n6553 = n2583 & n6552;
  assign n6554 = n100 & n6553;
  assign n6555 = ~n667 & n6554;
  assign n6556 = ~n641 & n6555;
  assign n6557 = ~n189 & n6556;
  assign n6558 = ~n107 & n6557;
  assign n6559 = ~n777 & n6558;
  assign n6560 = ~n564 & n6559;
  assign n6561 = ~n81 & n6560;
  assign n6562 = n423 & ~n1062;
  assign n6563 = ~n884 & n6562;
  assign n6564 = ~n298 & n6563;
  assign n6565 = ~n525 & n6564;
  assign n6566 = ~n284 & n1128;
  assign n6567 = ~n460 & n6566;
  assign n6568 = n1740 & n3416;
  assign n6569 = n2220 & n6568;
  assign n6570 = n6567 & n6569;
  assign n6571 = n1692 & n6570;
  assign n6572 = n6565 & n6571;
  assign n6573 = n877 & n6572;
  assign n6574 = n1709 & n6573;
  assign n6575 = n268 & n6574;
  assign n6576 = n4367 & n6575;
  assign n6577 = n6561 & n6576;
  assign n6578 = n5063 & n6577;
  assign n6579 = n450 & n6578;
  assign n6580 = n1761 & n6579;
  assign n6581 = ~n194 & n6580;
  assign n6582 = ~n151 & n6581;
  assign n6583 = ~n275 & n6582;
  assign n6584 = ~n173 & n6583;
  assign n6585 = ~n493 & n6584;
  assign n6586 = ~n200 & n6585;
  assign n6587 = ~n2388 & n3020;
  assign n6588 = ~n2464 & n3028;
  assign n6589 = ~n2533 & n3023;
  assign n6590 = n2844 & ~n2846;
  assign n6591 = ~n2847 & ~n6590;
  assign n6592 = n75 & n6591;
  assign n6593 = ~n6589 & ~n6592;
  assign n6594 = ~n6588 & n6593;
  assign n6595 = ~n6587 & n6594;
  assign n6596 = ~n6586 & ~n6595;
  assign n6597 = n918 & n2191;
  assign n6598 = n279 & n6597;
  assign n6599 = n100 & n6598;
  assign n6600 = ~n289 & n6599;
  assign n6601 = ~n803 & n6600;
  assign n6602 = ~n246 & n6601;
  assign n6603 = ~n466 & n6602;
  assign n6604 = ~n672 & n6603;
  assign n6605 = ~n328 & n515;
  assign n6606 = ~n396 & n6605;
  assign n6607 = ~n468 & n6606;
  assign n6608 = ~n752 & n1824;
  assign n6609 = ~n716 & n6608;
  assign n6610 = ~n489 & n6609;
  assign n6611 = n1424 & n1588;
  assign n6612 = n6610 & n6611;
  assign n6613 = n6607 & n6612;
  assign n6614 = n5148 & n6613;
  assign n6615 = n720 & n6614;
  assign n6616 = n634 & n6615;
  assign n6617 = ~n398 & n6616;
  assign n6618 = ~n152 & n6617;
  assign n6619 = ~n354 & n6618;
  assign n6620 = ~n777 & n6619;
  assign n6621 = ~n416 & n6620;
  assign n6622 = ~n368 & n6621;
  assign n6623 = ~n932 & n6622;
  assign n6624 = ~n272 & n6623;
  assign n6625 = ~n712 & n6624;
  assign n6626 = ~n558 & n2169;
  assign n6627 = ~n339 & n6626;
  assign n6628 = ~n327 & n6627;
  assign n6629 = n172 & n1497;
  assign n6630 = n6628 & n6629;
  assign n6631 = n2370 & n6630;
  assign n6632 = n3768 & n6631;
  assign n6633 = n5224 & n6632;
  assign n6634 = n6625 & n6633;
  assign n6635 = n6604 & n6634;
  assign n6636 = ~n353 & n6635;
  assign n6637 = ~n367 & n6636;
  assign n6638 = ~n825 & n6637;
  assign n6639 = ~n191 & n6638;
  assign n6640 = ~n225 & n6639;
  assign n6641 = ~n436 & n6640;
  assign n6642 = ~n2464 & n3020;
  assign n6643 = ~n2533 & n3028;
  assign n6644 = ~n2571 & n3023;
  assign n6645 = n2840 & ~n2842;
  assign n6646 = ~n2843 & ~n6645;
  assign n6647 = n75 & n6646;
  assign n6648 = ~n6644 & ~n6647;
  assign n6649 = ~n6643 & n6648;
  assign n6650 = ~n6642 & n6649;
  assign n6651 = ~n6641 & ~n6650;
  assign n6652 = n3314 & n3549;
  assign n6653 = n3409 & n6652;
  assign n6654 = n1105 & n6653;
  assign n6655 = n1523 & n6654;
  assign n6656 = ~n123 & n6655;
  assign n6657 = ~n427 & n6656;
  assign n6658 = ~n329 & n6657;
  assign n6659 = ~n328 & n6658;
  assign n6660 = ~n402 & n6659;
  assign n6661 = ~n430 & n6660;
  assign n6662 = ~n340 & n6661;
  assign n6663 = ~n358 & ~n518;
  assign n6664 = ~n428 & n6663;
  assign n6665 = n827 & n6664;
  assign n6666 = ~n306 & n6665;
  assign n6667 = ~n158 & n6666;
  assign n6668 = ~n161 & ~n531;
  assign n6669 = ~n304 & n6668;
  assign n6670 = ~n222 & n6669;
  assign n6671 = ~n280 & n604;
  assign n6672 = ~n332 & n6671;
  assign n6673 = n1578 & n6672;
  assign n6674 = n4269 & n6673;
  assign n6675 = n6670 & n6674;
  assign n6676 = n6667 & n6675;
  assign n6677 = n2258 & n6676;
  assign n6678 = n6662 & n6677;
  assign n6679 = n805 & n6678;
  assign n6680 = n2573 & n6679;
  assign n6681 = n1531 & n6680;
  assign n6682 = n1141 & n6681;
  assign n6683 = n978 & n6682;
  assign n6684 = n1161 & n6683;
  assign n6685 = ~n353 & n6684;
  assign n6686 = ~n299 & n6685;
  assign n6687 = ~n490 & n6686;
  assign n6688 = ~n568 & n6687;
  assign n6689 = ~n164 & n6688;
  assign n6690 = ~n623 & n6689;
  assign n6691 = ~n2533 & n3020;
  assign n6692 = ~n2571 & n3028;
  assign n6693 = ~n2674 & n3023;
  assign n6694 = n2836 & ~n2838;
  assign n6695 = ~n2839 & ~n6694;
  assign n6696 = n75 & n6695;
  assign n6697 = ~n6693 & ~n6696;
  assign n6698 = ~n6692 & n6697;
  assign n6699 = ~n6691 & n6698;
  assign n6700 = ~n6690 & ~n6699;
  assign n6701 = n300 & ~n301;
  assign n6702 = ~n1102 & n6701;
  assign n6703 = ~n203 & n6702;
  assign n6704 = ~n326 & n6703;
  assign n6705 = ~n287 & n6704;
  assign n6706 = ~n145 & ~n164;
  assign n6707 = ~n536 & n6706;
  assign n6708 = n1528 & n1617;
  assign n6709 = n2633 & n6708;
  assign n6710 = n3886 & n6709;
  assign n6711 = ~n715 & n6710;
  assign n6712 = ~n372 & n6711;
  assign n6713 = ~n366 & n6712;
  assign n6714 = ~n633 & n6713;
  assign n6715 = ~n132 & n3581;
  assign n6716 = ~n201 & n6715;
  assign n6717 = ~n557 & n2089;
  assign n6718 = n2423 & n6717;
  assign n6719 = n6716 & n6718;
  assign n6720 = n897 & n6719;
  assign n6721 = n1476 & n6720;
  assign n6722 = n665 & n6721;
  assign n6723 = n6714 & n6722;
  assign n6724 = n1531 & n6723;
  assign n6725 = n826 & n6724;
  assign n6726 = n227 & n6725;
  assign n6727 = ~n518 & n6726;
  assign n6728 = ~n1101 & n6727;
  assign n6729 = ~n192 & n6728;
  assign n6730 = ~n932 & n6729;
  assign n6731 = ~n474 & n6730;
  assign n6732 = ~n532 & n6731;
  assign n6733 = ~n233 & n885;
  assign n6734 = ~n144 & n6733;
  assign n6735 = n1221 & n6734;
  assign n6736 = n1615 & n6735;
  assign n6737 = n2632 & n6736;
  assign n6738 = n1454 & n6737;
  assign n6739 = n6732 & n6738;
  assign n6740 = n6707 & n6739;
  assign n6741 = n2021 & n6740;
  assign n6742 = n6705 & n6741;
  assign n6743 = ~n331 & n6742;
  assign n6744 = ~n272 & n6743;
  assign n6745 = ~n451 & n6744;
  assign n6746 = ~n1104 & n6745;
  assign n6747 = ~n562 & n6746;
  assign n6748 = ~n655 & n6747;
  assign n6749 = n300 & n2704;
  assign n6750 = ~n111 & n6749;
  assign n6751 = ~n1306 & n6750;
  assign n6752 = ~n374 & n6751;
  assign n6753 = ~n563 & n6752;
  assign n6754 = ~n331 & n6753;
  assign n6755 = ~n371 & n6754;
  assign n6756 = n5201 & n5793;
  assign n6757 = n776 & n6756;
  assign n6758 = n467 & n6757;
  assign n6759 = n6670 & n6758;
  assign n6760 = n2738 & n6759;
  assign n6761 = n873 & n6760;
  assign n6762 = n2010 & n6761;
  assign n6763 = n1824 & n6762;
  assign n6764 = n2073 & n6763;
  assign n6765 = ~n716 & n6764;
  assign n6766 = ~n422 & n6765;
  assign n6767 = ~n394 & n6766;
  assign n6768 = ~n603 & n6767;
  assign n6769 = ~n883 & n6768;
  assign n6770 = ~n1127 & n3636;
  assign n6771 = ~n633 & n6770;
  assign n6772 = n735 & n1586;
  assign n6773 = n6771 & n6772;
  assign n6774 = n4148 & n6773;
  assign n6775 = n2104 & n6774;
  assign n6776 = n6769 & n6775;
  assign n6777 = n6755 & n6776;
  assign n6778 = n510 & n6777;
  assign n6779 = n1668 & n6778;
  assign n6780 = n288 & n6779;
  assign n6781 = n869 & n6780;
  assign n6782 = n2466 & n6781;
  assign n6783 = n810 & n6782;
  assign n6784 = ~n236 & n6783;
  assign n6785 = ~n289 & n6784;
  assign n6786 = ~n254 & n6785;
  assign n6787 = ~n511 & n6786;
  assign n6788 = ~n203 & n6787;
  assign n6789 = ~n367 & n6788;
  assign n6790 = ~n777 & n6789;
  assign n6791 = ~n246 & n6790;
  assign n6792 = ~n2674 & n3020;
  assign n6793 = ~n2736 & n3028;
  assign n6794 = ~n2829 & n3023;
  assign n6795 = ~n2736 & n2829;
  assign n6796 = n2674 & ~n6795;
  assign n6797 = n2737 & n2829;
  assign n6798 = ~n6796 & ~n6797;
  assign n6799 = n75 & n6798;
  assign n6800 = ~n6794 & ~n6799;
  assign n6801 = ~n6793 & n6800;
  assign n6802 = ~n6792 & n6801;
  assign n6803 = ~n6791 & ~n6802;
  assign n6804 = ~n6748 & n6803;
  assign n6805 = n2832 & ~n2834;
  assign n6806 = ~n2835 & ~n6805;
  assign n6807 = n75 & n6806;
  assign n6808 = ~n2571 & n3020;
  assign n6809 = ~n2736 & n3023;
  assign n6810 = ~n2674 & n3028;
  assign n6811 = ~n6809 & ~n6810;
  assign n6812 = ~n6808 & n6811;
  assign n6813 = ~n6807 & n6812;
  assign n6814 = n6748 & ~n6803;
  assign n6815 = ~n6804 & ~n6814;
  assign n6816 = ~n6813 & n6815;
  assign n6817 = ~n6804 & ~n6816;
  assign n6818 = ~n6690 & ~n6700;
  assign n6819 = ~n6699 & ~n6700;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = ~n6817 & ~n6820;
  assign n6822 = ~n6700 & ~n6821;
  assign n6823 = ~n6641 & ~n6651;
  assign n6824 = ~n6650 & ~n6651;
  assign n6825 = ~n6823 & ~n6824;
  assign n6826 = ~n6822 & ~n6825;
  assign n6827 = ~n6651 & ~n6826;
  assign n6828 = ~n6586 & ~n6596;
  assign n6829 = ~n6595 & ~n6596;
  assign n6830 = ~n6828 & ~n6829;
  assign n6831 = ~n6827 & ~n6830;
  assign n6832 = ~n6596 & ~n6831;
  assign n6833 = ~n6536 & ~n6546;
  assign n6834 = ~n6545 & ~n6546;
  assign n6835 = ~n6833 & ~n6834;
  assign n6836 = ~n6832 & ~n6835;
  assign n6837 = ~n6546 & ~n6836;
  assign n6838 = ~n6500 & ~n6837;
  assign n6839 = n6500 & n6837;
  assign n6840 = ~n6838 & ~n6839;
  assign n6841 = ~n1992 & n3457;
  assign n6842 = ~n2152 & n3542;
  assign n6843 = ~n2057 & n3606;
  assign n6844 = ~n6842 & ~n6843;
  assign n6845 = ~n6841 & n6844;
  assign n6846 = ~n3368 & n6845;
  assign n6847 = ~n6143 & n6845;
  assign n6848 = ~n6846 & ~n6847;
  assign n6849 =  a[29]  & ~n6848;
  assign n6850 = ~ a[29]  & n6848;
  assign n6851 = ~n6849 & ~n6850;
  assign n6852 = n6840 & ~n6851;
  assign n6853 = ~n6838 & ~n6852;
  assign n6854 = ~n6487 & ~n6497;
  assign n6855 = ~n6496 & ~n6497;
  assign n6856 = ~n6854 & ~n6855;
  assign n6857 = ~n6853 & ~n6856;
  assign n6858 = ~n6497 & ~n6857;
  assign n6859 = ~n6474 & ~n6484;
  assign n6860 = ~n6483 & ~n6484;
  assign n6861 = ~n6859 & ~n6860;
  assign n6862 = ~n6858 & ~n6861;
  assign n6863 = ~n6484 & ~n6862;
  assign n6864 = ~n6471 & ~n6863;
  assign n6865 = n6471 & n6863;
  assign n6866 = ~n6864 & ~n6865;
  assign n6867 = ~n1779 & n3457;
  assign n6868 = ~n1913 & n3542;
  assign n6869 = ~n1877 & n3606;
  assign n6870 = ~n6868 & ~n6869;
  assign n6871 = ~n6867 & n6870;
  assign n6872 = n3368 & n5851;
  assign n6873 = n6871 & ~n6872;
  assign n6874 =  a[29]  & ~n6873;
  assign n6875 =  a[29]  & ~n6874;
  assign n6876 = ~n6873 & ~n6874;
  assign n6877 = ~n6875 & ~n6876;
  assign n6878 = n6866 & ~n6877;
  assign n6879 = ~n6864 & ~n6878;
  assign n6880 = ~n6157 & n6168;
  assign n6881 = ~n6169 & ~n6880;
  assign n6882 = ~n6879 & n6881;
  assign n6883 = n6879 & ~n6881;
  assign n6884 = ~n6882 & ~n6883;
  assign n6885 = ~n1364 & n3884;
  assign n6886 = ~n1572 & n3967;
  assign n6887 = ~n1472 & n4046;
  assign n6888 = ~n6886 & ~n6887;
  assign n6889 = ~n6885 & n6888;
  assign n6890 = n4050 & n5114;
  assign n6891 = n6889 & ~n6890;
  assign n6892 =  a[26]  & ~n6891;
  assign n6893 =  a[26]  & ~n6892;
  assign n6894 = ~n6891 & ~n6892;
  assign n6895 = ~n6893 & ~n6894;
  assign n6896 = n6884 & ~n6895;
  assign n6897 = ~n6882 & ~n6896;
  assign n6898 = ~n6468 & ~n6897;
  assign n6899 = n6468 & n6897;
  assign n6900 = ~n6898 & ~n6899;
  assign n6901 = ~n958 & n4694;
  assign n6902 = ~n1178 & n4533;
  assign n6903 = ~n1060 & n4604;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = ~n6901 & n6904;
  assign n6906 = n4536 & n4633;
  assign n6907 = n6905 & ~n6906;
  assign n6908 =  a[23]  & ~n6907;
  assign n6909 =  a[23]  & ~n6908;
  assign n6910 = ~n6907 & ~n6908;
  assign n6911 = ~n6909 & ~n6910;
  assign n6912 = n6900 & ~n6911;
  assign n6913 = ~n6898 & ~n6912;
  assign n6914 = ~n6465 & ~n6913;
  assign n6915 = ~n6462 & ~n6914;
  assign n6916 = ~n6448 & ~n6915;
  assign n6917 = n6448 & n6915;
  assign n6918 = ~n6916 & ~n6917;
  assign n6919 = ~n3012 & n5496;
  assign n6920 = ~n587 & n4935;
  assign n6921 = ~n392 & n5407;
  assign n6922 = ~n6920 & ~n6921;
  assign n6923 = ~n6919 & n6922;
  assign n6924 = n3018 & n4938;
  assign n6925 = n6923 & ~n6924;
  assign n6926 =  a[20]  & ~n6925;
  assign n6927 =  a[20]  & ~n6926;
  assign n6928 = ~n6925 & ~n6926;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = n6918 & ~n6929;
  assign n6931 = ~n6916 & ~n6930;
  assign n6932 = ~n6445 & ~n6931;
  assign n6933 = n6445 & n6931;
  assign n6934 = ~n6932 & ~n6933;
  assign n6935 = ~n3805 & n6233;
  assign n6936 = ~n3605 & n5663;
  assign n6937 = ~n3456 & n5939;
  assign n6938 = ~n6936 & ~n6937;
  assign n6939 = ~n6935 & n6938;
  assign n6940 = n3818 & n5666;
  assign n6941 = n6939 & ~n6940;
  assign n6942 =  a[17]  & ~n6941;
  assign n6943 =  a[17]  & ~n6942;
  assign n6944 = ~n6941 & ~n6942;
  assign n6945 = ~n6943 & ~n6944;
  assign n6946 = n6934 & ~n6945;
  assign n6947 = ~n6932 & ~n6946;
  assign n6948 = ~n6442 & ~n6947;
  assign n6949 = ~n6439 & ~n6948;
  assign n6950 = ~n3877 & n6402;
  assign n6951 = n6393 & ~n6400;
  assign n6952 = ~n4515 & n6951;
  assign n6953 = ~n6950 & ~n6952;
  assign n6954 = ~n6397 & n6953;
  assign n6955 = ~n4609 & n6953;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 =  a[14]  & ~n6956;
  assign n6958 = ~ a[14]  & n6956;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = ~n6949 & ~n6959;
  assign n6961 = n6377 & ~n6389;
  assign n6962 = ~n6388 & ~n6389;
  assign n6963 = ~n6961 & ~n6962;
  assign n6964 = n6949 & n6959;
  assign n6965 = ~n6960 & ~n6964;
  assign n6966 = ~n6963 & n6965;
  assign n6967 = ~n6960 & ~n6966;
  assign n6968 = ~n6425 & ~n6967;
  assign n6969 = n6425 & n6967;
  assign n6970 = ~n6968 & ~n6969;
  assign n6971 = n6934 & ~n6946;
  assign n6972 = ~n6945 & ~n6946;
  assign n6973 = ~n6971 & ~n6972;
  assign n6974 = n6918 & ~n6930;
  assign n6975 = ~n6929 & ~n6930;
  assign n6976 = ~n6974 & ~n6975;
  assign n6977 = n6465 & n6913;
  assign n6978 = ~n6914 & ~n6977;
  assign n6979 = ~n392 & n5496;
  assign n6980 = ~n710 & n4935;
  assign n6981 = ~n587 & n5407;
  assign n6982 = ~n6980 & ~n6981;
  assign n6983 = ~n6979 & n6982;
  assign n6984 = ~n4938 & n6983;
  assign n6985 = ~n3347 & n6983;
  assign n6986 = ~n6984 & ~n6985;
  assign n6987 =  a[20]  & ~n6986;
  assign n6988 = ~ a[20]  & n6986;
  assign n6989 = ~n6987 & ~n6988;
  assign n6990 = n6978 & ~n6989;
  assign n6991 = n6900 & ~n6912;
  assign n6992 = ~n6911 & ~n6912;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = n6884 & ~n6896;
  assign n6995 = ~n6895 & ~n6896;
  assign n6996 = ~n6994 & ~n6995;
  assign n6997 = n6866 & ~n6878;
  assign n6998 = ~n6877 & ~n6878;
  assign n6999 = ~n6997 & ~n6998;
  assign n7000 = ~n1472 & n3884;
  assign n7001 = ~n1665 & n3967;
  assign n7002 = ~n1572 & n4046;
  assign n7003 = ~n7001 & ~n7002;
  assign n7004 = ~n7000 & n7003;
  assign n7005 = ~n4050 & n7004;
  assign n7006 = ~n5139 & n7004;
  assign n7007 = ~n7005 & ~n7006;
  assign n7008 =  a[26]  & ~n7007;
  assign n7009 = ~ a[26]  & n7007;
  assign n7010 = ~n7008 & ~n7009;
  assign n7011 = ~n6999 & ~n7010;
  assign n7012 = ~n6858 & ~n6862;
  assign n7013 = ~n6861 & ~n6862;
  assign n7014 = ~n7012 & ~n7013;
  assign n7015 = ~n1877 & n3457;
  assign n7016 = ~n1992 & n3542;
  assign n7017 = ~n1913 & n3606;
  assign n7018 = ~n7016 & ~n7017;
  assign n7019 = ~n7015 & n7018;
  assign n7020 = ~n3368 & n7019;
  assign n7021 = ~n6007 & n7019;
  assign n7022 = ~n7020 & ~n7021;
  assign n7023 =  a[29]  & ~n7022;
  assign n7024 = ~ a[29]  & n7022;
  assign n7025 = ~n7023 & ~n7024;
  assign n7026 = ~n7014 & ~n7025;
  assign n7027 = n7014 & n7025;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = ~n1572 & n3884;
  assign n7030 = ~n1779 & n3967;
  assign n7031 = ~n1665 & n4046;
  assign n7032 = ~n7030 & ~n7031;
  assign n7033 = ~n7029 & n7032;
  assign n7034 = n4050 & n5561;
  assign n7035 = n7033 & ~n7034;
  assign n7036 =  a[26]  & ~n7035;
  assign n7037 =  a[26]  & ~n7036;
  assign n7038 = ~n7035 & ~n7036;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = n7028 & ~n7039;
  assign n7041 = ~n7026 & ~n7040;
  assign n7042 = n6999 & n7010;
  assign n7043 = ~n7011 & ~n7042;
  assign n7044 = ~n7041 & n7043;
  assign n7045 = ~n7011 & ~n7044;
  assign n7046 = ~n6996 & ~n7045;
  assign n7047 = n6996 & n7045;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = ~n1060 & n4694;
  assign n7050 = ~n1235 & n4533;
  assign n7051 = ~n1178 & n4604;
  assign n7052 = ~n7050 & ~n7051;
  assign n7053 = ~n7049 & n7052;
  assign n7054 = n4429 & n4536;
  assign n7055 = n7053 & ~n7054;
  assign n7056 =  a[23]  & ~n7055;
  assign n7057 =  a[23]  & ~n7056;
  assign n7058 = ~n7055 & ~n7056;
  assign n7059 = ~n7057 & ~n7058;
  assign n7060 = n7048 & ~n7059;
  assign n7061 = ~n7046 & ~n7060;
  assign n7062 = ~n6993 & ~n7061;
  assign n7063 = n6993 & n7061;
  assign n7064 = ~n7062 & ~n7063;
  assign n7065 = ~n587 & n5496;
  assign n7066 = ~n867 & n4935;
  assign n7067 = ~n710 & n5407;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = ~n7065 & n7068;
  assign n7070 = n3331 & n4938;
  assign n7071 = n7069 & ~n7070;
  assign n7072 =  a[20]  & ~n7071;
  assign n7073 =  a[20]  & ~n7072;
  assign n7074 = ~n7071 & ~n7072;
  assign n7075 = ~n7073 & ~n7074;
  assign n7076 = n7064 & ~n7075;
  assign n7077 = ~n7062 & ~n7076;
  assign n7078 = ~n6978 & n6989;
  assign n7079 = ~n6990 & ~n7078;
  assign n7080 = ~n7077 & n7079;
  assign n7081 = ~n6990 & ~n7080;
  assign n7082 = ~n6976 & ~n7081;
  assign n7083 = n6976 & n7081;
  assign n7084 = ~n7082 & ~n7083;
  assign n7085 = ~n3456 & n6233;
  assign n7086 = ~n3539 & n5663;
  assign n7087 = ~n3605 & n5939;
  assign n7088 = ~n7086 & ~n7087;
  assign n7089 = ~n7085 & n7088;
  assign n7090 = n3627 & n5666;
  assign n7091 = n7089 & ~n7090;
  assign n7092 =  a[17]  & ~n7091;
  assign n7093 =  a[17]  & ~n7092;
  assign n7094 = ~n7091 & ~n7092;
  assign n7095 = ~n7093 & ~n7094;
  assign n7096 = n7084 & ~n7095;
  assign n7097 = ~n7082 & ~n7096;
  assign n7098 = ~n6973 & ~n7097;
  assign n7099 = n6973 & n7097;
  assign n7100 = ~n7098 & ~n7099;
  assign n7101 = ~n6393 & n6396;
  assign n7102 = ~n3877 & n7101;
  assign n7103 = ~n3964 & n6402;
  assign n7104 = ~n4045 & n6951;
  assign n7105 = ~n7103 & ~n7104;
  assign n7106 = ~n7102 & n7105;
  assign n7107 = n4067 & n6397;
  assign n7108 = n7106 & ~n7107;
  assign n7109 =  a[14]  & ~n7108;
  assign n7110 =  a[14]  & ~n7109;
  assign n7111 = ~n7108 & ~n7109;
  assign n7112 = ~n7110 & ~n7111;
  assign n7113 = n7100 & ~n7112;
  assign n7114 = ~n7098 & ~n7113;
  assign n7115 = ~n4515 & n7101;
  assign n7116 = ~n4045 & n6402;
  assign n7117 = ~n3877 & n6951;
  assign n7118 = ~n7116 & ~n7117;
  assign n7119 = ~n7115 & n7118;
  assign n7120 = ~n6397 & n7119;
  assign n7121 = ~n4715 & n7119;
  assign n7122 = ~n7120 & ~n7121;
  assign n7123 =  a[14]  & ~n7122;
  assign n7124 = ~ a[14]  & n7122;
  assign n7125 = ~n7123 & ~n7124;
  assign n7126 = ~n7114 & ~n7125;
  assign n7127 = n6442 & n6947;
  assign n7128 = ~n6948 & ~n7127;
  assign n7129 = ~n7114 & ~n7126;
  assign n7130 = ~n7125 & ~n7126;
  assign n7131 = ~n7129 & ~n7130;
  assign n7132 = n7128 & ~n7131;
  assign n7133 = ~n7126 & ~n7132;
  assign n7134 = n6963 & ~n6965;
  assign n7135 = ~n6966 & ~n7134;
  assign n7136 = ~n7133 & n7135;
  assign n7137 = n7084 & ~n7096;
  assign n7138 = ~n7095 & ~n7096;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = ~n3605 & n6233;
  assign n7141 = ~n3012 & n5663;
  assign n7142 = ~n3539 & n5939;
  assign n7143 = ~n7141 & ~n7142;
  assign n7144 = ~n7140 & n7143;
  assign n7145 = n4084 & n5666;
  assign n7146 = n7144 & ~n7145;
  assign n7147 =  a[17]  & ~n7146;
  assign n7148 = ~n7146 & ~n7147;
  assign n7149 =  a[17]  & ~n7147;
  assign n7150 = ~n7148 & ~n7149;
  assign n7151 = n7077 & ~n7079;
  assign n7152 = ~n7080 & ~n7151;
  assign n7153 = ~n7150 & n7152;
  assign n7154 = ~n7150 & ~n7153;
  assign n7155 = n7152 & ~n7153;
  assign n7156 = ~n7154 & ~n7155;
  assign n7157 = n7064 & ~n7076;
  assign n7158 = ~n7075 & ~n7076;
  assign n7159 = ~n7157 & ~n7158;
  assign n7160 = n7048 & ~n7060;
  assign n7161 = ~n7059 & ~n7060;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~n1178 & n4694;
  assign n7164 = ~n1364 & n4533;
  assign n7165 = ~n1235 & n4604;
  assign n7166 = ~n7164 & ~n7165;
  assign n7167 = ~n7163 & n7166;
  assign n7168 = n4536 & n4861;
  assign n7169 = n7167 & ~n7168;
  assign n7170 =  a[23]  & ~n7169;
  assign n7171 = ~n7169 & ~n7170;
  assign n7172 =  a[23]  & ~n7170;
  assign n7173 = ~n7171 & ~n7172;
  assign n7174 = n7041 & ~n7043;
  assign n7175 = ~n7044 & ~n7174;
  assign n7176 = ~n7173 & n7175;
  assign n7177 = ~n7173 & ~n7176;
  assign n7178 = n7175 & ~n7176;
  assign n7179 = ~n7177 & ~n7178;
  assign n7180 = n7028 & ~n7040;
  assign n7181 = ~n7039 & ~n7040;
  assign n7182 = ~n7180 & ~n7181;
  assign n7183 = ~n6853 & ~n6857;
  assign n7184 = ~n6856 & ~n6857;
  assign n7185 = ~n7183 & ~n7184;
  assign n7186 = ~n1913 & n3457;
  assign n7187 = ~n2057 & n3542;
  assign n7188 = ~n1992 & n3606;
  assign n7189 = ~n7187 & ~n7188;
  assign n7190 = ~n7186 & n7189;
  assign n7191 = ~n3368 & n7190;
  assign n7192 = ~n5834 & n7190;
  assign n7193 = ~n7191 & ~n7192;
  assign n7194 =  a[29]  & ~n7193;
  assign n7195 = ~ a[29]  & n7193;
  assign n7196 = ~n7194 & ~n7195;
  assign n7197 = ~n7185 & ~n7196;
  assign n7198 = n7185 & n7196;
  assign n7199 = ~n7197 & ~n7198;
  assign n7200 = ~n1665 & n3884;
  assign n7201 = ~n1877 & n3967;
  assign n7202 = ~n1779 & n4046;
  assign n7203 = ~n7201 & ~n7202;
  assign n7204 = ~n7200 & n7203;
  assign n7205 = n4050 & n5328;
  assign n7206 = n7204 & ~n7205;
  assign n7207 =  a[26]  & ~n7206;
  assign n7208 =  a[26]  & ~n7207;
  assign n7209 = ~n7206 & ~n7207;
  assign n7210 = ~n7208 & ~n7209;
  assign n7211 = n7199 & ~n7210;
  assign n7212 = ~n7197 & ~n7211;
  assign n7213 = ~n7182 & ~n7212;
  assign n7214 = n7182 & n7212;
  assign n7215 = ~n7213 & ~n7214;
  assign n7216 = ~n1235 & n4694;
  assign n7217 = ~n1472 & n4533;
  assign n7218 = ~n1364 & n4604;
  assign n7219 = ~n7217 & ~n7218;
  assign n7220 = ~n7216 & n7219;
  assign n7221 = n4536 & n4848;
  assign n7222 = n7220 & ~n7221;
  assign n7223 =  a[23]  & ~n7222;
  assign n7224 =  a[23]  & ~n7223;
  assign n7225 = ~n7222 & ~n7223;
  assign n7226 = ~n7224 & ~n7225;
  assign n7227 = n7215 & ~n7226;
  assign n7228 = ~n7213 & ~n7227;
  assign n7229 = ~n7179 & ~n7228;
  assign n7230 = ~n7176 & ~n7229;
  assign n7231 = ~n7162 & ~n7230;
  assign n7232 = n7162 & n7230;
  assign n7233 = ~n7231 & ~n7232;
  assign n7234 = ~n710 & n5496;
  assign n7235 = ~n958 & n4935;
  assign n7236 = ~n867 & n5407;
  assign n7237 = ~n7235 & ~n7236;
  assign n7238 = ~n7234 & n7237;
  assign n7239 = n4179 & n4938;
  assign n7240 = n7238 & ~n7239;
  assign n7241 =  a[20]  & ~n7240;
  assign n7242 =  a[20]  & ~n7241;
  assign n7243 = ~n7240 & ~n7241;
  assign n7244 = ~n7242 & ~n7243;
  assign n7245 = n7233 & ~n7244;
  assign n7246 = ~n7231 & ~n7245;
  assign n7247 = ~n7159 & ~n7246;
  assign n7248 = n7159 & n7246;
  assign n7249 = ~n7247 & ~n7248;
  assign n7250 = ~n3539 & n6233;
  assign n7251 = ~n392 & n5663;
  assign n7252 = ~n3012 & n5939;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = ~n7250 & n7253;
  assign n7255 = n3715 & n5666;
  assign n7256 = n7254 & ~n7255;
  assign n7257 =  a[17]  & ~n7256;
  assign n7258 =  a[17]  & ~n7257;
  assign n7259 = ~n7256 & ~n7257;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = n7249 & ~n7260;
  assign n7262 = ~n7247 & ~n7261;
  assign n7263 = ~n7156 & ~n7262;
  assign n7264 = ~n7153 & ~n7263;
  assign n7265 = ~n7139 & ~n7264;
  assign n7266 = n7139 & n7264;
  assign n7267 = ~n7265 & ~n7266;
  assign n7268 = ~n4045 & n7101;
  assign n7269 = ~n3805 & n6402;
  assign n7270 = ~n3964 & n6951;
  assign n7271 = ~n7269 & ~n7270;
  assign n7272 = ~n7268 & n7271;
  assign n7273 = n4477 & n6397;
  assign n7274 = n7272 & ~n7273;
  assign n7275 =  a[14]  & ~n7274;
  assign n7276 =  a[14]  & ~n7275;
  assign n7277 = ~n7274 & ~n7275;
  assign n7278 = ~n7276 & ~n7277;
  assign n7279 = n7267 & ~n7278;
  assign n7280 = ~n7265 & ~n7279;
  assign n7281 = ~ a[9]  &  a[10] ;
  assign n7282 =  a[9]  & ~ a[10] ;
  assign n7283 = ~n7281 & ~n7282;
  assign n7284 =  a[10]  & ~ a[11] ;
  assign n7285 = ~ a[10]  &  a[11] ;
  assign n7286 = ~n7284 & ~n7285;
  assign n7287 =  a[8]  & ~ a[9] ;
  assign n7288 = ~ a[8]  &  a[9] ;
  assign n7289 = ~n7287 & ~n7288;
  assign n7290 = ~n7286 & n7289;
  assign n7291 = n7283 & n7290;
  assign n7292 = ~n4515 & n7291;
  assign n7293 = ~n4522 & ~n7292;
  assign n7294 = ~n7286 & ~n7289;
  assign n7295 = ~n7292 & ~n7294;
  assign n7296 = ~n7293 & ~n7295;
  assign n7297 =  a[11]  & ~n7296;
  assign n7298 = ~ a[11]  & n7296;
  assign n7299 = ~n7297 & ~n7298;
  assign n7300 = ~n7280 & ~n7299;
  assign n7301 = n7100 & ~n7113;
  assign n7302 = ~n7112 & ~n7113;
  assign n7303 = ~n7301 & ~n7302;
  assign n7304 = n7280 & n7299;
  assign n7305 = ~n7300 & ~n7304;
  assign n7306 = ~n7303 & n7305;
  assign n7307 = ~n7300 & ~n7306;
  assign n7308 = ~n7128 & ~n7130;
  assign n7309 = ~n7129 & n7308;
  assign n7310 = ~n7132 & ~n7309;
  assign n7311 = ~n7307 & n7310;
  assign n7312 = ~n7303 & ~n7306;
  assign n7313 = n7305 & ~n7306;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = n7156 & n7262;
  assign n7316 = ~n7263 & ~n7315;
  assign n7317 = ~n3964 & n7101;
  assign n7318 = ~n3456 & n6402;
  assign n7319 = ~n3805 & n6951;
  assign n7320 = ~n7318 & ~n7319;
  assign n7321 = ~n7317 & n7320;
  assign n7322 = ~n6397 & n7321;
  assign n7323 = ~n4558 & n7321;
  assign n7324 = ~n7322 & ~n7323;
  assign n7325 =  a[14]  & ~n7324;
  assign n7326 = ~ a[14]  & n7324;
  assign n7327 = ~n7325 & ~n7326;
  assign n7328 = n7316 & ~n7327;
  assign n7329 = n7249 & ~n7261;
  assign n7330 = ~n7260 & ~n7261;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = n7233 & ~n7245;
  assign n7333 = ~n7244 & ~n7245;
  assign n7334 = ~n7332 & ~n7333;
  assign n7335 = n7179 & n7228;
  assign n7336 = ~n7229 & ~n7335;
  assign n7337 = ~n867 & n5496;
  assign n7338 = ~n1060 & n4935;
  assign n7339 = ~n958 & n5407;
  assign n7340 = ~n7338 & ~n7339;
  assign n7341 = ~n7337 & n7340;
  assign n7342 = ~n4938 & n7341;
  assign n7343 = ~n4204 & n7341;
  assign n7344 = ~n7342 & ~n7343;
  assign n7345 =  a[20]  & ~n7344;
  assign n7346 = ~ a[20]  & n7344;
  assign n7347 = ~n7345 & ~n7346;
  assign n7348 = n7336 & ~n7347;
  assign n7349 = n7215 & ~n7227;
  assign n7350 = ~n7226 & ~n7227;
  assign n7351 = ~n7349 & ~n7350;
  assign n7352 = n7199 & ~n7211;
  assign n7353 = ~n7210 & ~n7211;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = ~n6832 & ~n6836;
  assign n7356 = ~n6835 & ~n6836;
  assign n7357 = ~n7355 & ~n7356;
  assign n7358 = ~n2057 & n3457;
  assign n7359 = ~n2189 & n3542;
  assign n7360 = ~n2152 & n3606;
  assign n7361 = ~n7359 & ~n7360;
  assign n7362 = ~n7358 & n7361;
  assign n7363 = ~n3368 & n7362;
  assign n7364 = ~n6479 & n7362;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 =  a[29]  & ~n7365;
  assign n7367 = ~ a[29]  & n7365;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = ~n7357 & ~n7368;
  assign n7370 = ~n6827 & ~n6831;
  assign n7371 = ~n6830 & ~n6831;
  assign n7372 = ~n7370 & ~n7371;
  assign n7373 = ~n2152 & n3457;
  assign n7374 = ~n2291 & n3542;
  assign n7375 = ~n2189 & n3606;
  assign n7376 = ~n7374 & ~n7375;
  assign n7377 = ~n7373 & n7376;
  assign n7378 = ~n3368 & n7377;
  assign n7379 = ~n6492 & n7377;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 =  a[29]  & ~n7380;
  assign n7382 = ~ a[29]  & n7380;
  assign n7383 = ~n7381 & ~n7382;
  assign n7384 = ~n7372 & ~n7383;
  assign n7385 = ~n2189 & n3457;
  assign n7386 = ~n2388 & n3542;
  assign n7387 = ~n2291 & n3606;
  assign n7388 = ~n7386 & ~n7387;
  assign n7389 = ~n7385 & n7388;
  assign n7390 = n3368 & n6122;
  assign n7391 = n7389 & ~n7390;
  assign n7392 =  a[29]  & ~n7391;
  assign n7393 = ~n7391 & ~n7392;
  assign n7394 =  a[29]  & ~n7392;
  assign n7395 = ~n7393 & ~n7394;
  assign n7396 = ~n6822 & ~n6826;
  assign n7397 = ~n6825 & ~n6826;
  assign n7398 = ~n7396 & ~n7397;
  assign n7399 = ~n7395 & ~n7398;
  assign n7400 = ~n7395 & ~n7399;
  assign n7401 = ~n7398 & ~n7399;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = ~n2291 & n3457;
  assign n7404 = ~n2464 & n3542;
  assign n7405 = ~n2388 & n3606;
  assign n7406 = ~n7404 & ~n7405;
  assign n7407 = ~n7403 & n7406;
  assign n7408 = n3368 & n6541;
  assign n7409 = n7407 & ~n7408;
  assign n7410 =  a[29]  & ~n7409;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 =  a[29]  & ~n7410;
  assign n7413 = ~n7411 & ~n7412;
  assign n7414 = ~n6817 & ~n6821;
  assign n7415 = ~n6820 & ~n6821;
  assign n7416 = ~n7414 & ~n7415;
  assign n7417 = ~n7413 & ~n7416;
  assign n7418 = ~n7413 & ~n7417;
  assign n7419 = ~n7416 & ~n7417;
  assign n7420 = ~n7418 & ~n7419;
  assign n7421 = ~n2388 & n3457;
  assign n7422 = ~n2533 & n3542;
  assign n7423 = ~n2464 & n3606;
  assign n7424 = ~n7422 & ~n7423;
  assign n7425 = ~n7421 & n7424;
  assign n7426 = n3368 & n6591;
  assign n7427 = n7425 & ~n7426;
  assign n7428 =  a[29]  & ~n7427;
  assign n7429 = ~n7427 & ~n7428;
  assign n7430 =  a[29]  & ~n7428;
  assign n7431 = ~n7429 & ~n7430;
  assign n7432 = ~n6813 & ~n6816;
  assign n7433 = n6815 & ~n6816;
  assign n7434 = ~n7432 & ~n7433;
  assign n7435 = ~n7431 & ~n7434;
  assign n7436 = ~n7431 & ~n7435;
  assign n7437 = ~n7434 & ~n7435;
  assign n7438 = ~n7436 & ~n7437;
  assign n7439 = ~n2464 & n3457;
  assign n7440 = ~n2571 & n3542;
  assign n7441 = ~n2533 & n3606;
  assign n7442 = ~n7440 & ~n7441;
  assign n7443 = ~n7439 & n7442;
  assign n7444 = n3368 & n6646;
  assign n7445 = n7443 & ~n7444;
  assign n7446 =  a[29]  & ~n7445;
  assign n7447 = ~n7445 & ~n7446;
  assign n7448 =  a[29]  & ~n7446;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = ~n6791 & ~n6803;
  assign n7451 = ~n6802 & ~n6803;
  assign n7452 = ~n7450 & ~n7451;
  assign n7453 = ~n7449 & ~n7452;
  assign n7454 = ~n7449 & ~n7453;
  assign n7455 = ~n7452 & ~n7453;
  assign n7456 = ~n7454 & ~n7455;
  assign n7457 = ~n2533 & n3457;
  assign n7458 = ~n2674 & n3542;
  assign n7459 = ~n2571 & n3606;
  assign n7460 = ~n7458 & ~n7459;
  assign n7461 = ~n7457 & n7460;
  assign n7462 = n3368 & n6695;
  assign n7463 = n7461 & ~n7462;
  assign n7464 =  a[29]  & ~n7463;
  assign n7465 = ~n7463 & ~n7464;
  assign n7466 =  a[29]  & ~n7464;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = n2736 & ~n2829;
  assign n7469 = ~n6795 & ~n7468;
  assign n7470 = n75 & ~n7469;
  assign n7471 = ~n2829 & n3028;
  assign n7472 = ~n2736 & n3020;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = ~n7470 & n7473;
  assign n7475 = ~n7467 & ~n7474;
  assign n7476 = ~n7467 & ~n7475;
  assign n7477 = ~n7474 & ~n7475;
  assign n7478 = ~n7476 & ~n7477;
  assign n7479 = ~n75 & ~n3020;
  assign n7480 = ~n2829 & ~n7479;
  assign n7481 = ~n2829 & n3606;
  assign n7482 = ~n2736 & n3457;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = n3368 & ~n7469;
  assign n7485 = n7483 & ~n7484;
  assign n7486 =  a[29]  & ~n7485;
  assign n7487 =  a[29]  & ~n7486;
  assign n7488 = ~n7485 & ~n7486;
  assign n7489 = ~n7487 & ~n7488;
  assign n7490 = ~n2829 & ~n3367;
  assign n7491 =  a[29]  & ~n7490;
  assign n7492 = ~n7489 & n7491;
  assign n7493 = ~n2674 & n3457;
  assign n7494 = ~n2829 & n3542;
  assign n7495 = ~n2736 & n3606;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n7493 & n7496;
  assign n7498 = ~n3368 & n7497;
  assign n7499 = ~n6798 & n7497;
  assign n7500 = ~n7498 & ~n7499;
  assign n7501 =  a[29]  & ~n7500;
  assign n7502 = ~ a[29]  & n7500;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = n7492 & ~n7503;
  assign n7505 = n7480 & n7504;
  assign n7506 = ~n2571 & n3457;
  assign n7507 = ~n2736 & n3542;
  assign n7508 = ~n2674 & n3606;
  assign n7509 = ~n7507 & ~n7508;
  assign n7510 = ~n7506 & n7509;
  assign n7511 = n3368 & n6806;
  assign n7512 = n7510 & ~n7511;
  assign n7513 =  a[29]  & ~n7512;
  assign n7514 = ~n7512 & ~n7513;
  assign n7515 =  a[29]  & ~n7513;
  assign n7516 = ~n7514 & ~n7515;
  assign n7517 = ~n7480 & n7504;
  assign n7518 = n7480 & ~n7504;
  assign n7519 = ~n7517 & ~n7518;
  assign n7520 = ~n7516 & ~n7519;
  assign n7521 = ~n7505 & ~n7520;
  assign n7522 = ~n7478 & ~n7521;
  assign n7523 = ~n7475 & ~n7522;
  assign n7524 = ~n7456 & ~n7523;
  assign n7525 = ~n7453 & ~n7524;
  assign n7526 = ~n7438 & ~n7525;
  assign n7527 = ~n7435 & ~n7526;
  assign n7528 = ~n7420 & ~n7527;
  assign n7529 = ~n7417 & ~n7528;
  assign n7530 = ~n7402 & ~n7529;
  assign n7531 = ~n7399 & ~n7530;
  assign n7532 = n7372 & n7383;
  assign n7533 = ~n7384 & ~n7532;
  assign n7534 = ~n7531 & n7533;
  assign n7535 = ~n7384 & ~n7534;
  assign n7536 = n7357 & n7368;
  assign n7537 = ~n7369 & ~n7536;
  assign n7538 = ~n7535 & n7537;
  assign n7539 = ~n7369 & ~n7538;
  assign n7540 = ~n6840 & n6851;
  assign n7541 = ~n6852 & ~n7540;
  assign n7542 = ~n7539 & n7541;
  assign n7543 = ~n1779 & n3884;
  assign n7544 = ~n1913 & n3967;
  assign n7545 = ~n1877 & n4046;
  assign n7546 = ~n7544 & ~n7545;
  assign n7547 = ~n7543 & n7546;
  assign n7548 = n4050 & n5851;
  assign n7549 = n7547 & ~n7548;
  assign n7550 =  a[26]  & ~n7549;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 =  a[26]  & ~n7550;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = n7539 & ~n7541;
  assign n7555 = ~n7542 & ~n7554;
  assign n7556 = ~n7553 & n7555;
  assign n7557 = ~n7542 & ~n7556;
  assign n7558 = ~n7354 & ~n7557;
  assign n7559 = n7354 & n7557;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = ~n1364 & n4694;
  assign n7562 = ~n1572 & n4533;
  assign n7563 = ~n1472 & n4604;
  assign n7564 = ~n7562 & ~n7563;
  assign n7565 = ~n7561 & n7564;
  assign n7566 = n4536 & n5114;
  assign n7567 = n7565 & ~n7566;
  assign n7568 =  a[23]  & ~n7567;
  assign n7569 =  a[23]  & ~n7568;
  assign n7570 = ~n7567 & ~n7568;
  assign n7571 = ~n7569 & ~n7570;
  assign n7572 = n7560 & ~n7571;
  assign n7573 = ~n7558 & ~n7572;
  assign n7574 = ~n7351 & ~n7573;
  assign n7575 = n7351 & n7573;
  assign n7576 = ~n7574 & ~n7575;
  assign n7577 = ~n958 & n5496;
  assign n7578 = ~n1178 & n4935;
  assign n7579 = ~n1060 & n5407;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = ~n7577 & n7580;
  assign n7582 = n4633 & n4938;
  assign n7583 = n7581 & ~n7582;
  assign n7584 =  a[20]  & ~n7583;
  assign n7585 =  a[20]  & ~n7584;
  assign n7586 = ~n7583 & ~n7584;
  assign n7587 = ~n7585 & ~n7586;
  assign n7588 = n7576 & ~n7587;
  assign n7589 = ~n7574 & ~n7588;
  assign n7590 = ~n7336 & n7347;
  assign n7591 = ~n7348 & ~n7590;
  assign n7592 = ~n7589 & n7591;
  assign n7593 = ~n7348 & ~n7592;
  assign n7594 = ~n7334 & ~n7593;
  assign n7595 = n7334 & n7593;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~n3012 & n6233;
  assign n7598 = ~n587 & n5663;
  assign n7599 = ~n392 & n5939;
  assign n7600 = ~n7598 & ~n7599;
  assign n7601 = ~n7597 & n7600;
  assign n7602 = n3018 & n5666;
  assign n7603 = n7601 & ~n7602;
  assign n7604 =  a[17]  & ~n7603;
  assign n7605 =  a[17]  & ~n7604;
  assign n7606 = ~n7603 & ~n7604;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = n7596 & ~n7607;
  assign n7609 = ~n7594 & ~n7608;
  assign n7610 = ~n7331 & ~n7609;
  assign n7611 = n7331 & n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~n3805 & n7101;
  assign n7614 = ~n3605 & n6402;
  assign n7615 = ~n3456 & n6951;
  assign n7616 = ~n7614 & ~n7615;
  assign n7617 = ~n7613 & n7616;
  assign n7618 = n3818 & n6397;
  assign n7619 = n7617 & ~n7618;
  assign n7620 =  a[14]  & ~n7619;
  assign n7621 =  a[14]  & ~n7620;
  assign n7622 = ~n7619 & ~n7620;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = n7612 & ~n7623;
  assign n7625 = ~n7610 & ~n7624;
  assign n7626 = n7316 & ~n7328;
  assign n7627 = ~n7327 & ~n7328;
  assign n7628 = ~n7626 & ~n7627;
  assign n7629 = ~n7625 & ~n7628;
  assign n7630 = ~n7328 & ~n7629;
  assign n7631 = ~n3877 & n7291;
  assign n7632 = ~n7283 & n7289;
  assign n7633 = ~n4515 & n7632;
  assign n7634 = ~n7631 & ~n7633;
  assign n7635 = ~n7294 & n7634;
  assign n7636 = ~n4609 & n7634;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 =  a[11]  & ~n7637;
  assign n7639 = ~ a[11]  & n7637;
  assign n7640 = ~n7638 & ~n7639;
  assign n7641 = ~n7630 & ~n7640;
  assign n7642 = n7267 & ~n7279;
  assign n7643 = ~n7278 & ~n7279;
  assign n7644 = ~n7642 & ~n7643;
  assign n7645 = n7630 & n7640;
  assign n7646 = ~n7641 & ~n7645;
  assign n7647 = ~n7644 & n7646;
  assign n7648 = ~n7641 & ~n7647;
  assign n7649 = ~n7314 & ~n7648;
  assign n7650 = n7314 & n7648;
  assign n7651 = ~n7649 & ~n7650;
  assign n7652 = n7612 & ~n7624;
  assign n7653 = ~n7623 & ~n7624;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = n7596 & ~n7608;
  assign n7656 = ~n7607 & ~n7608;
  assign n7657 = ~n7655 & ~n7656;
  assign n7658 = ~n392 & n6233;
  assign n7659 = ~n710 & n5663;
  assign n7660 = ~n587 & n5939;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n7658 & n7661;
  assign n7663 = n3347 & n5666;
  assign n7664 = n7662 & ~n7663;
  assign n7665 =  a[17]  & ~n7664;
  assign n7666 = ~n7664 & ~n7665;
  assign n7667 =  a[17]  & ~n7665;
  assign n7668 = ~n7666 & ~n7667;
  assign n7669 = n7589 & ~n7591;
  assign n7670 = ~n7592 & ~n7669;
  assign n7671 = ~n7668 & n7670;
  assign n7672 = ~n7668 & ~n7671;
  assign n7673 = n7670 & ~n7671;
  assign n7674 = ~n7672 & ~n7673;
  assign n7675 = n7576 & ~n7588;
  assign n7676 = ~n7587 & ~n7588;
  assign n7677 = ~n7675 & ~n7676;
  assign n7678 = n7560 & ~n7572;
  assign n7679 = ~n7571 & ~n7572;
  assign n7680 = ~n7678 & ~n7679;
  assign n7681 = n7535 & ~n7537;
  assign n7682 = ~n7538 & ~n7681;
  assign n7683 = ~n1877 & n3884;
  assign n7684 = ~n1992 & n3967;
  assign n7685 = ~n1913 & n4046;
  assign n7686 = ~n7684 & ~n7685;
  assign n7687 = ~n7683 & n7686;
  assign n7688 = ~n4050 & n7687;
  assign n7689 = ~n6007 & n7687;
  assign n7690 = ~n7688 & ~n7689;
  assign n7691 =  a[26]  & ~n7690;
  assign n7692 = ~ a[26]  & n7690;
  assign n7693 = ~n7691 & ~n7692;
  assign n7694 = n7682 & ~n7693;
  assign n7695 = n7531 & ~n7533;
  assign n7696 = ~n7534 & ~n7695;
  assign n7697 = ~n1913 & n3884;
  assign n7698 = ~n2057 & n3967;
  assign n7699 = ~n1992 & n4046;
  assign n7700 = ~n7698 & ~n7699;
  assign n7701 = ~n7697 & n7700;
  assign n7702 = ~n4050 & n7701;
  assign n7703 = ~n5834 & n7701;
  assign n7704 = ~n7702 & ~n7703;
  assign n7705 =  a[26]  & ~n7704;
  assign n7706 = ~ a[26]  & n7704;
  assign n7707 = ~n7705 & ~n7706;
  assign n7708 = n7696 & ~n7707;
  assign n7709 = n7402 & n7529;
  assign n7710 = ~n7530 & ~n7709;
  assign n7711 = ~n1992 & n3884;
  assign n7712 = ~n2152 & n3967;
  assign n7713 = ~n2057 & n4046;
  assign n7714 = ~n7712 & ~n7713;
  assign n7715 = ~n7711 & n7714;
  assign n7716 = ~n4050 & n7715;
  assign n7717 = ~n6143 & n7715;
  assign n7718 = ~n7716 & ~n7717;
  assign n7719 =  a[26]  & ~n7718;
  assign n7720 = ~ a[26]  & n7718;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = n7710 & ~n7721;
  assign n7723 = n7420 & n7527;
  assign n7724 = ~n7528 & ~n7723;
  assign n7725 = ~n2057 & n3884;
  assign n7726 = ~n2189 & n3967;
  assign n7727 = ~n2152 & n4046;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = ~n7725 & n7728;
  assign n7730 = ~n4050 & n7729;
  assign n7731 = ~n6479 & n7729;
  assign n7732 = ~n7730 & ~n7731;
  assign n7733 =  a[26]  & ~n7732;
  assign n7734 = ~ a[26]  & n7732;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = n7724 & ~n7735;
  assign n7737 = n7438 & n7525;
  assign n7738 = ~n7526 & ~n7737;
  assign n7739 = ~n2152 & n3884;
  assign n7740 = ~n2291 & n3967;
  assign n7741 = ~n2189 & n4046;
  assign n7742 = ~n7740 & ~n7741;
  assign n7743 = ~n7739 & n7742;
  assign n7744 = ~n4050 & n7743;
  assign n7745 = ~n6492 & n7743;
  assign n7746 = ~n7744 & ~n7745;
  assign n7747 =  a[26]  & ~n7746;
  assign n7748 = ~ a[26]  & n7746;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = n7738 & ~n7749;
  assign n7751 = n7456 & n7523;
  assign n7752 = ~n7524 & ~n7751;
  assign n7753 = ~n2189 & n3884;
  assign n7754 = ~n2388 & n3967;
  assign n7755 = ~n2291 & n4046;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = ~n7753 & n7756;
  assign n7758 = ~n4050 & n7757;
  assign n7759 = ~n6122 & n7757;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 =  a[26]  & ~n7760;
  assign n7762 = ~ a[26]  & n7760;
  assign n7763 = ~n7761 & ~n7762;
  assign n7764 = n7752 & ~n7763;
  assign n7765 = ~n7478 & ~n7522;
  assign n7766 = ~n7521 & ~n7522;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = ~n2291 & n3884;
  assign n7769 = ~n2464 & n3967;
  assign n7770 = ~n2388 & n4046;
  assign n7771 = ~n7769 & ~n7770;
  assign n7772 = ~n7768 & n7771;
  assign n7773 = ~n4050 & n7772;
  assign n7774 = ~n6541 & n7772;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 =  a[26]  & ~n7775;
  assign n7777 = ~ a[26]  & n7775;
  assign n7778 = ~n7776 & ~n7777;
  assign n7779 = ~n7767 & ~n7778;
  assign n7780 = ~n2388 & n3884;
  assign n7781 = ~n2533 & n3967;
  assign n7782 = ~n2464 & n4046;
  assign n7783 = ~n7781 & ~n7782;
  assign n7784 = ~n7780 & n7783;
  assign n7785 = n4050 & n6591;
  assign n7786 = n7784 & ~n7785;
  assign n7787 =  a[26]  & ~n7786;
  assign n7788 = ~n7786 & ~n7787;
  assign n7789 =  a[26]  & ~n7787;
  assign n7790 = ~n7788 & ~n7789;
  assign n7791 = n7516 & n7519;
  assign n7792 = ~n7520 & ~n7791;
  assign n7793 = ~n7790 & n7792;
  assign n7794 = ~n7790 & ~n7793;
  assign n7795 = n7792 & ~n7793;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = ~n2464 & n3884;
  assign n7798 = ~n2571 & n3967;
  assign n7799 = ~n2533 & n4046;
  assign n7800 = ~n7798 & ~n7799;
  assign n7801 = ~n7797 & n7800;
  assign n7802 = n4050 & n6646;
  assign n7803 = n7801 & ~n7802;
  assign n7804 =  a[26]  & ~n7803;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 =  a[26]  & ~n7804;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = ~n7492 & n7503;
  assign n7809 = ~n7504 & ~n7808;
  assign n7810 = ~n7807 & n7809;
  assign n7811 = ~n7807 & ~n7810;
  assign n7812 = n7809 & ~n7810;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = n7489 & ~n7491;
  assign n7815 = ~n7492 & ~n7814;
  assign n7816 = ~n2533 & n3884;
  assign n7817 = ~n2674 & n3967;
  assign n7818 = ~n2571 & n4046;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = ~n7816 & n7819;
  assign n7821 = ~n4050 & n7820;
  assign n7822 = ~n6695 & n7820;
  assign n7823 = ~n7821 & ~n7822;
  assign n7824 =  a[26]  & ~n7823;
  assign n7825 = ~ a[26]  & n7823;
  assign n7826 = ~n7824 & ~n7825;
  assign n7827 = n7815 & ~n7826;
  assign n7828 = ~n2829 & n4046;
  assign n7829 = ~n2736 & n3884;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = n4050 & ~n7469;
  assign n7832 = n7830 & ~n7831;
  assign n7833 =  a[26]  & ~n7832;
  assign n7834 =  a[26]  & ~n7833;
  assign n7835 = ~n7832 & ~n7833;
  assign n7836 = ~n7834 & ~n7835;
  assign n7837 = ~n2829 & ~n3880;
  assign n7838 =  a[26]  & ~n7837;
  assign n7839 = ~n7836 & n7838;
  assign n7840 = ~n2674 & n3884;
  assign n7841 = ~n2829 & n3967;
  assign n7842 = ~n2736 & n4046;
  assign n7843 = ~n7841 & ~n7842;
  assign n7844 = ~n7840 & n7843;
  assign n7845 = ~n4050 & n7844;
  assign n7846 = ~n6798 & n7844;
  assign n7847 = ~n7845 & ~n7846;
  assign n7848 =  a[26]  & ~n7847;
  assign n7849 = ~ a[26]  & n7847;
  assign n7850 = ~n7848 & ~n7849;
  assign n7851 = n7839 & ~n7850;
  assign n7852 = n7490 & n7851;
  assign n7853 = n7851 & ~n7852;
  assign n7854 = n7490 & ~n7852;
  assign n7855 = ~n7853 & ~n7854;
  assign n7856 = ~n2571 & n3884;
  assign n7857 = ~n2736 & n3967;
  assign n7858 = ~n2674 & n4046;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n7856 & n7859;
  assign n7861 = n4050 & n6806;
  assign n7862 = n7860 & ~n7861;
  assign n7863 =  a[26]  & ~n7862;
  assign n7864 =  a[26]  & ~n7863;
  assign n7865 = ~n7862 & ~n7863;
  assign n7866 = ~n7864 & ~n7865;
  assign n7867 = ~n7855 & ~n7866;
  assign n7868 = ~n7852 & ~n7867;
  assign n7869 = ~n7815 & n7826;
  assign n7870 = ~n7827 & ~n7869;
  assign n7871 = ~n7868 & n7870;
  assign n7872 = ~n7827 & ~n7871;
  assign n7873 = ~n7813 & ~n7872;
  assign n7874 = ~n7810 & ~n7873;
  assign n7875 = ~n7796 & ~n7874;
  assign n7876 = ~n7793 & ~n7875;
  assign n7877 = ~n7767 & ~n7779;
  assign n7878 = ~n7778 & ~n7779;
  assign n7879 = ~n7877 & ~n7878;
  assign n7880 = ~n7876 & ~n7879;
  assign n7881 = ~n7779 & ~n7880;
  assign n7882 = n7752 & ~n7764;
  assign n7883 = ~n7763 & ~n7764;
  assign n7884 = ~n7882 & ~n7883;
  assign n7885 = ~n7881 & ~n7884;
  assign n7886 = ~n7764 & ~n7885;
  assign n7887 = n7738 & ~n7750;
  assign n7888 = ~n7749 & ~n7750;
  assign n7889 = ~n7887 & ~n7888;
  assign n7890 = ~n7886 & ~n7889;
  assign n7891 = ~n7750 & ~n7890;
  assign n7892 = n7724 & ~n7736;
  assign n7893 = ~n7735 & ~n7736;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = ~n7891 & ~n7894;
  assign n7896 = ~n7736 & ~n7895;
  assign n7897 = n7710 & ~n7722;
  assign n7898 = ~n7721 & ~n7722;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = ~n7896 & ~n7899;
  assign n7901 = ~n7722 & ~n7900;
  assign n7902 = n7696 & ~n7708;
  assign n7903 = ~n7707 & ~n7708;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = ~n7901 & ~n7904;
  assign n7906 = ~n7708 & ~n7905;
  assign n7907 = n7682 & ~n7694;
  assign n7908 = ~n7693 & ~n7694;
  assign n7909 = ~n7907 & ~n7908;
  assign n7910 = ~n7906 & ~n7909;
  assign n7911 = ~n7694 & ~n7910;
  assign n7912 = n7553 & ~n7555;
  assign n7913 = ~n7556 & ~n7912;
  assign n7914 = ~n7911 & n7913;
  assign n7915 = ~n1472 & n4694;
  assign n7916 = ~n1665 & n4533;
  assign n7917 = ~n1572 & n4604;
  assign n7918 = ~n7916 & ~n7917;
  assign n7919 = ~n7915 & n7918;
  assign n7920 = n4536 & n5139;
  assign n7921 = n7919 & ~n7920;
  assign n7922 =  a[23]  & ~n7921;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 =  a[23]  & ~n7922;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = n7911 & ~n7913;
  assign n7927 = ~n7914 & ~n7926;
  assign n7928 = ~n7925 & n7927;
  assign n7929 = ~n7914 & ~n7928;
  assign n7930 = ~n7680 & ~n7929;
  assign n7931 = n7680 & n7929;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = ~n1060 & n5496;
  assign n7934 = ~n1235 & n4935;
  assign n7935 = ~n1178 & n5407;
  assign n7936 = ~n7934 & ~n7935;
  assign n7937 = ~n7933 & n7936;
  assign n7938 = n4429 & n4938;
  assign n7939 = n7937 & ~n7938;
  assign n7940 =  a[20]  & ~n7939;
  assign n7941 =  a[20]  & ~n7940;
  assign n7942 = ~n7939 & ~n7940;
  assign n7943 = ~n7941 & ~n7942;
  assign n7944 = n7932 & ~n7943;
  assign n7945 = ~n7930 & ~n7944;
  assign n7946 = ~n7677 & ~n7945;
  assign n7947 = n7677 & n7945;
  assign n7948 = ~n7946 & ~n7947;
  assign n7949 = ~n587 & n6233;
  assign n7950 = ~n867 & n5663;
  assign n7951 = ~n710 & n5939;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = ~n7949 & n7952;
  assign n7954 = n3331 & n5666;
  assign n7955 = n7953 & ~n7954;
  assign n7956 =  a[17]  & ~n7955;
  assign n7957 =  a[17]  & ~n7956;
  assign n7958 = ~n7955 & ~n7956;
  assign n7959 = ~n7957 & ~n7958;
  assign n7960 = n7948 & ~n7959;
  assign n7961 = ~n7946 & ~n7960;
  assign n7962 = ~n7674 & ~n7961;
  assign n7963 = ~n7671 & ~n7962;
  assign n7964 = ~n7657 & ~n7963;
  assign n7965 = n7657 & n7963;
  assign n7966 = ~n7964 & ~n7965;
  assign n7967 = ~n3456 & n7101;
  assign n7968 = ~n3539 & n6402;
  assign n7969 = ~n3605 & n6951;
  assign n7970 = ~n7968 & ~n7969;
  assign n7971 = ~n7967 & n7970;
  assign n7972 = n3627 & n6397;
  assign n7973 = n7971 & ~n7972;
  assign n7974 =  a[14]  & ~n7973;
  assign n7975 =  a[14]  & ~n7974;
  assign n7976 = ~n7973 & ~n7974;
  assign n7977 = ~n7975 & ~n7976;
  assign n7978 = n7966 & ~n7977;
  assign n7979 = ~n7964 & ~n7978;
  assign n7980 = ~n7654 & ~n7979;
  assign n7981 = n7654 & n7979;
  assign n7982 = ~n7980 & ~n7981;
  assign n7983 = n7286 & ~n7289;
  assign n7984 = ~n3877 & n7983;
  assign n7985 = ~n3964 & n7291;
  assign n7986 = ~n4045 & n7632;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = ~n7984 & n7987;
  assign n7989 = n4067 & n7294;
  assign n7990 = n7988 & ~n7989;
  assign n7991 =  a[11]  & ~n7990;
  assign n7992 =  a[11]  & ~n7991;
  assign n7993 = ~n7990 & ~n7991;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = n7982 & ~n7994;
  assign n7996 = ~n7980 & ~n7995;
  assign n7997 = ~n4515 & n7983;
  assign n7998 = ~n4045 & n7291;
  assign n7999 = ~n3877 & n7632;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = ~n7997 & n8000;
  assign n8002 = ~n7294 & n8001;
  assign n8003 = ~n4715 & n8001;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 =  a[11]  & ~n8004;
  assign n8006 = ~ a[11]  & n8004;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = ~n7996 & ~n8007;
  assign n8009 = n7996 & n8007;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = ~n7625 & ~n7629;
  assign n8012 = ~n7628 & ~n7629;
  assign n8013 = ~n8011 & ~n8012;
  assign n8014 = n8010 & ~n8013;
  assign n8015 = ~n8008 & ~n8014;
  assign n8016 = n7644 & ~n7646;
  assign n8017 = ~n7647 & ~n8016;
  assign n8018 = ~n8015 & n8017;
  assign n8019 = n8010 & ~n8014;
  assign n8020 = ~n8013 & ~n8014;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = n7966 & ~n7978;
  assign n8023 = ~n7977 & ~n7978;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = n7674 & n7961;
  assign n8026 = ~n7962 & ~n8025;
  assign n8027 = ~n3605 & n7101;
  assign n8028 = ~n3012 & n6402;
  assign n8029 = ~n3539 & n6951;
  assign n8030 = ~n8028 & ~n8029;
  assign n8031 = ~n8027 & n8030;
  assign n8032 = ~n6397 & n8031;
  assign n8033 = ~n4084 & n8031;
  assign n8034 = ~n8032 & ~n8033;
  assign n8035 =  a[14]  & ~n8034;
  assign n8036 = ~ a[14]  & n8034;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = n8026 & ~n8037;
  assign n8039 = n7948 & ~n7960;
  assign n8040 = ~n7959 & ~n7960;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = n7932 & ~n7944;
  assign n8043 = ~n7943 & ~n7944;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = ~n1572 & n4694;
  assign n8046 = ~n1779 & n4533;
  assign n8047 = ~n1665 & n4604;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = ~n8045 & n8048;
  assign n8050 = n4536 & n5561;
  assign n8051 = n8049 & ~n8050;
  assign n8052 =  a[23]  & ~n8051;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 =  a[23]  & ~n8052;
  assign n8055 = ~n8053 & ~n8054;
  assign n8056 = ~n7906 & ~n7910;
  assign n8057 = ~n7909 & ~n7910;
  assign n8058 = ~n8056 & ~n8057;
  assign n8059 = ~n8055 & ~n8058;
  assign n8060 = ~n8055 & ~n8059;
  assign n8061 = ~n8058 & ~n8059;
  assign n8062 = ~n8060 & ~n8061;
  assign n8063 = ~n1665 & n4694;
  assign n8064 = ~n1877 & n4533;
  assign n8065 = ~n1779 & n4604;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = ~n8063 & n8066;
  assign n8068 = n4536 & n5328;
  assign n8069 = n8067 & ~n8068;
  assign n8070 =  a[23]  & ~n8069;
  assign n8071 = ~n8069 & ~n8070;
  assign n8072 =  a[23]  & ~n8070;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = ~n7901 & ~n7905;
  assign n8075 = ~n7904 & ~n7905;
  assign n8076 = ~n8074 & ~n8075;
  assign n8077 = ~n8073 & ~n8076;
  assign n8078 = ~n8073 & ~n8077;
  assign n8079 = ~n8076 & ~n8077;
  assign n8080 = ~n8078 & ~n8079;
  assign n8081 = ~n1779 & n4694;
  assign n8082 = ~n1913 & n4533;
  assign n8083 = ~n1877 & n4604;
  assign n8084 = ~n8082 & ~n8083;
  assign n8085 = ~n8081 & n8084;
  assign n8086 = n4536 & n5851;
  assign n8087 = n8085 & ~n8086;
  assign n8088 =  a[23]  & ~n8087;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 =  a[23]  & ~n8088;
  assign n8091 = ~n8089 & ~n8090;
  assign n8092 = ~n7896 & ~n7900;
  assign n8093 = ~n7899 & ~n7900;
  assign n8094 = ~n8092 & ~n8093;
  assign n8095 = ~n8091 & ~n8094;
  assign n8096 = ~n8091 & ~n8095;
  assign n8097 = ~n8094 & ~n8095;
  assign n8098 = ~n8096 & ~n8097;
  assign n8099 = ~n1877 & n4694;
  assign n8100 = ~n1992 & n4533;
  assign n8101 = ~n1913 & n4604;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = ~n8099 & n8102;
  assign n8104 = n4536 & n6007;
  assign n8105 = n8103 & ~n8104;
  assign n8106 =  a[23]  & ~n8105;
  assign n8107 = ~n8105 & ~n8106;
  assign n8108 =  a[23]  & ~n8106;
  assign n8109 = ~n8107 & ~n8108;
  assign n8110 = ~n7891 & ~n7895;
  assign n8111 = ~n7894 & ~n7895;
  assign n8112 = ~n8110 & ~n8111;
  assign n8113 = ~n8109 & ~n8112;
  assign n8114 = ~n8109 & ~n8113;
  assign n8115 = ~n8112 & ~n8113;
  assign n8116 = ~n8114 & ~n8115;
  assign n8117 = ~n1913 & n4694;
  assign n8118 = ~n2057 & n4533;
  assign n8119 = ~n1992 & n4604;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = ~n8117 & n8120;
  assign n8122 = n4536 & n5834;
  assign n8123 = n8121 & ~n8122;
  assign n8124 =  a[23]  & ~n8123;
  assign n8125 = ~n8123 & ~n8124;
  assign n8126 =  a[23]  & ~n8124;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = ~n7886 & ~n7890;
  assign n8129 = ~n7889 & ~n7890;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = ~n8127 & ~n8130;
  assign n8132 = ~n8127 & ~n8131;
  assign n8133 = ~n8130 & ~n8131;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = ~n1992 & n4694;
  assign n8136 = ~n2152 & n4533;
  assign n8137 = ~n2057 & n4604;
  assign n8138 = ~n8136 & ~n8137;
  assign n8139 = ~n8135 & n8138;
  assign n8140 = n4536 & n6143;
  assign n8141 = n8139 & ~n8140;
  assign n8142 =  a[23]  & ~n8141;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 =  a[23]  & ~n8142;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = ~n7881 & ~n7885;
  assign n8147 = ~n7884 & ~n7885;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = ~n8145 & ~n8148;
  assign n8150 = ~n8145 & ~n8149;
  assign n8151 = ~n8148 & ~n8149;
  assign n8152 = ~n8150 & ~n8151;
  assign n8153 = ~n2057 & n4694;
  assign n8154 = ~n2189 & n4533;
  assign n8155 = ~n2152 & n4604;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = ~n8153 & n8156;
  assign n8158 = n4536 & n6479;
  assign n8159 = n8157 & ~n8158;
  assign n8160 =  a[23]  & ~n8159;
  assign n8161 = ~n8159 & ~n8160;
  assign n8162 =  a[23]  & ~n8160;
  assign n8163 = ~n8161 & ~n8162;
  assign n8164 = ~n7876 & ~n7880;
  assign n8165 = ~n7879 & ~n7880;
  assign n8166 = ~n8164 & ~n8165;
  assign n8167 = ~n8163 & ~n8166;
  assign n8168 = ~n8163 & ~n8167;
  assign n8169 = ~n8166 & ~n8167;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = n7796 & n7874;
  assign n8172 = ~n7875 & ~n8171;
  assign n8173 = ~n2152 & n4694;
  assign n8174 = ~n2291 & n4533;
  assign n8175 = ~n2189 & n4604;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = ~n8173 & n8176;
  assign n8178 = ~n4536 & n8177;
  assign n8179 = ~n6492 & n8177;
  assign n8180 = ~n8178 & ~n8179;
  assign n8181 =  a[23]  & ~n8180;
  assign n8182 = ~ a[23]  & n8180;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = n8172 & ~n8183;
  assign n8185 = n7813 & n7872;
  assign n8186 = ~n7873 & ~n8185;
  assign n8187 = ~n2189 & n4694;
  assign n8188 = ~n2388 & n4533;
  assign n8189 = ~n2291 & n4604;
  assign n8190 = ~n8188 & ~n8189;
  assign n8191 = ~n8187 & n8190;
  assign n8192 = ~n4536 & n8191;
  assign n8193 = ~n6122 & n8191;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 =  a[23]  & ~n8194;
  assign n8196 = ~ a[23]  & n8194;
  assign n8197 = ~n8195 & ~n8196;
  assign n8198 = n8186 & ~n8197;
  assign n8199 = ~n2291 & n4694;
  assign n8200 = ~n2464 & n4533;
  assign n8201 = ~n2388 & n4604;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = ~n8199 & n8202;
  assign n8204 = n4536 & n6541;
  assign n8205 = n8203 & ~n8204;
  assign n8206 =  a[23]  & ~n8205;
  assign n8207 = ~n8205 & ~n8206;
  assign n8208 =  a[23]  & ~n8206;
  assign n8209 = ~n8207 & ~n8208;
  assign n8210 = n7868 & ~n7870;
  assign n8211 = ~n7871 & ~n8210;
  assign n8212 = ~n8209 & n8211;
  assign n8213 = ~n8209 & ~n8212;
  assign n8214 = n8211 & ~n8212;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = ~n7855 & ~n7867;
  assign n8217 = ~n7866 & ~n7867;
  assign n8218 = ~n8216 & ~n8217;
  assign n8219 = ~n2388 & n4694;
  assign n8220 = ~n2533 & n4533;
  assign n8221 = ~n2464 & n4604;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = ~n8219 & n8222;
  assign n8224 = ~n4536 & n8223;
  assign n8225 = ~n6591 & n8223;
  assign n8226 = ~n8224 & ~n8225;
  assign n8227 =  a[23]  & ~n8226;
  assign n8228 = ~ a[23]  & n8226;
  assign n8229 = ~n8227 & ~n8228;
  assign n8230 = ~n8218 & ~n8229;
  assign n8231 = ~n2464 & n4694;
  assign n8232 = ~n2571 & n4533;
  assign n8233 = ~n2533 & n4604;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = ~n8231 & n8234;
  assign n8236 = n4536 & n6646;
  assign n8237 = n8235 & ~n8236;
  assign n8238 =  a[23]  & ~n8237;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 =  a[23]  & ~n8238;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = ~n7839 & n7850;
  assign n8243 = ~n7851 & ~n8242;
  assign n8244 = ~n8241 & n8243;
  assign n8245 = ~n8241 & ~n8244;
  assign n8246 = n8243 & ~n8244;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = n7836 & ~n7838;
  assign n8249 = ~n7839 & ~n8248;
  assign n8250 = ~n2533 & n4694;
  assign n8251 = ~n2674 & n4533;
  assign n8252 = ~n2571 & n4604;
  assign n8253 = ~n8251 & ~n8252;
  assign n8254 = ~n8250 & n8253;
  assign n8255 = ~n4536 & n8254;
  assign n8256 = ~n6695 & n8254;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 =  a[23]  & ~n8257;
  assign n8259 = ~ a[23]  & n8257;
  assign n8260 = ~n8258 & ~n8259;
  assign n8261 = n8249 & ~n8260;
  assign n8262 = ~n2829 & n4604;
  assign n8263 = ~n2736 & n4694;
  assign n8264 = ~n8262 & ~n8263;
  assign n8265 = n4536 & ~n7469;
  assign n8266 = n8264 & ~n8265;
  assign n8267 =  a[23]  & ~n8266;
  assign n8268 =  a[23]  & ~n8267;
  assign n8269 = ~n8266 & ~n8267;
  assign n8270 = ~n8268 & ~n8269;
  assign n8271 = ~n2829 & ~n4528;
  assign n8272 =  a[23]  & ~n8271;
  assign n8273 = ~n8270 & n8272;
  assign n8274 = ~n2674 & n4694;
  assign n8275 = ~n2829 & n4533;
  assign n8276 = ~n2736 & n4604;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = ~n8274 & n8277;
  assign n8279 = ~n4536 & n8278;
  assign n8280 = ~n6798 & n8278;
  assign n8281 = ~n8279 & ~n8280;
  assign n8282 =  a[23]  & ~n8281;
  assign n8283 = ~ a[23]  & n8281;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = n8273 & ~n8284;
  assign n8286 = n7837 & n8285;
  assign n8287 = n8285 & ~n8286;
  assign n8288 = n7837 & ~n8286;
  assign n8289 = ~n8287 & ~n8288;
  assign n8290 = ~n2571 & n4694;
  assign n8291 = ~n2736 & n4533;
  assign n8292 = ~n2674 & n4604;
  assign n8293 = ~n8291 & ~n8292;
  assign n8294 = ~n8290 & n8293;
  assign n8295 = n4536 & n6806;
  assign n8296 = n8294 & ~n8295;
  assign n8297 =  a[23]  & ~n8296;
  assign n8298 =  a[23]  & ~n8297;
  assign n8299 = ~n8296 & ~n8297;
  assign n8300 = ~n8298 & ~n8299;
  assign n8301 = ~n8289 & ~n8300;
  assign n8302 = ~n8286 & ~n8301;
  assign n8303 = ~n8249 & n8260;
  assign n8304 = ~n8261 & ~n8303;
  assign n8305 = ~n8302 & n8304;
  assign n8306 = ~n8261 & ~n8305;
  assign n8307 = ~n8247 & ~n8306;
  assign n8308 = ~n8244 & ~n8307;
  assign n8309 = n8218 & n8229;
  assign n8310 = ~n8230 & ~n8309;
  assign n8311 = ~n8308 & n8310;
  assign n8312 = ~n8230 & ~n8311;
  assign n8313 = ~n8215 & ~n8312;
  assign n8314 = ~n8212 & ~n8313;
  assign n8315 = n8186 & ~n8198;
  assign n8316 = ~n8197 & ~n8198;
  assign n8317 = ~n8315 & ~n8316;
  assign n8318 = ~n8314 & ~n8317;
  assign n8319 = ~n8198 & ~n8318;
  assign n8320 = ~n8172 & n8183;
  assign n8321 = ~n8184 & ~n8320;
  assign n8322 = ~n8319 & n8321;
  assign n8323 = ~n8184 & ~n8322;
  assign n8324 = ~n8170 & ~n8323;
  assign n8325 = ~n8167 & ~n8324;
  assign n8326 = ~n8152 & ~n8325;
  assign n8327 = ~n8149 & ~n8326;
  assign n8328 = ~n8134 & ~n8327;
  assign n8329 = ~n8131 & ~n8328;
  assign n8330 = ~n8116 & ~n8329;
  assign n8331 = ~n8113 & ~n8330;
  assign n8332 = ~n8098 & ~n8331;
  assign n8333 = ~n8095 & ~n8332;
  assign n8334 = ~n8080 & ~n8333;
  assign n8335 = ~n8077 & ~n8334;
  assign n8336 = ~n8062 & ~n8335;
  assign n8337 = ~n8059 & ~n8336;
  assign n8338 = n7925 & ~n7927;
  assign n8339 = ~n7928 & ~n8338;
  assign n8340 = ~n8337 & n8339;
  assign n8341 = ~n1178 & n5496;
  assign n8342 = ~n1364 & n4935;
  assign n8343 = ~n1235 & n5407;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = ~n8341 & n8344;
  assign n8346 = n4861 & n4938;
  assign n8347 = n8345 & ~n8346;
  assign n8348 =  a[20]  & ~n8347;
  assign n8349 = ~n8347 & ~n8348;
  assign n8350 =  a[20]  & ~n8348;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = n8337 & ~n8339;
  assign n8353 = ~n8340 & ~n8352;
  assign n8354 = ~n8351 & n8353;
  assign n8355 = ~n8340 & ~n8354;
  assign n8356 = ~n8044 & ~n8355;
  assign n8357 = n8044 & n8355;
  assign n8358 = ~n8356 & ~n8357;
  assign n8359 = ~n710 & n6233;
  assign n8360 = ~n958 & n5663;
  assign n8361 = ~n867 & n5939;
  assign n8362 = ~n8360 & ~n8361;
  assign n8363 = ~n8359 & n8362;
  assign n8364 = n4179 & n5666;
  assign n8365 = n8363 & ~n8364;
  assign n8366 =  a[17]  & ~n8365;
  assign n8367 =  a[17]  & ~n8366;
  assign n8368 = ~n8365 & ~n8366;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = n8358 & ~n8369;
  assign n8371 = ~n8356 & ~n8370;
  assign n8372 = ~n8041 & ~n8371;
  assign n8373 = n8041 & n8371;
  assign n8374 = ~n8372 & ~n8373;
  assign n8375 = ~n3539 & n7101;
  assign n8376 = ~n392 & n6402;
  assign n8377 = ~n3012 & n6951;
  assign n8378 = ~n8376 & ~n8377;
  assign n8379 = ~n8375 & n8378;
  assign n8380 = n3715 & n6397;
  assign n8381 = n8379 & ~n8380;
  assign n8382 =  a[14]  & ~n8381;
  assign n8383 =  a[14]  & ~n8382;
  assign n8384 = ~n8381 & ~n8382;
  assign n8385 = ~n8383 & ~n8384;
  assign n8386 = n8374 & ~n8385;
  assign n8387 = ~n8372 & ~n8386;
  assign n8388 = ~n8026 & n8037;
  assign n8389 = ~n8038 & ~n8388;
  assign n8390 = ~n8387 & n8389;
  assign n8391 = ~n8038 & ~n8390;
  assign n8392 = ~n8024 & ~n8391;
  assign n8393 = n8024 & n8391;
  assign n8394 = ~n8392 & ~n8393;
  assign n8395 = ~n4045 & n7983;
  assign n8396 = ~n3805 & n7291;
  assign n8397 = ~n3964 & n7632;
  assign n8398 = ~n8396 & ~n8397;
  assign n8399 = ~n8395 & n8398;
  assign n8400 = n4477 & n7294;
  assign n8401 = n8399 & ~n8400;
  assign n8402 =  a[11]  & ~n8401;
  assign n8403 =  a[11]  & ~n8402;
  assign n8404 = ~n8401 & ~n8402;
  assign n8405 = ~n8403 & ~n8404;
  assign n8406 = n8394 & ~n8405;
  assign n8407 = ~n8392 & ~n8406;
  assign n8408 = ~ a[6]  &  a[7] ;
  assign n8409 =  a[6]  & ~ a[7] ;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 =  a[7]  & ~ a[8] ;
  assign n8412 = ~ a[7]  &  a[8] ;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 =  a[5]  & ~ a[6] ;
  assign n8415 = ~ a[5]  &  a[6] ;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = ~n8413 & n8416;
  assign n8418 = n8410 & n8417;
  assign n8419 = ~n4515 & n8418;
  assign n8420 = ~n4522 & ~n8419;
  assign n8421 = ~n8413 & ~n8416;
  assign n8422 = ~n8419 & ~n8421;
  assign n8423 = ~n8420 & ~n8422;
  assign n8424 =  a[8]  & ~n8423;
  assign n8425 = ~ a[8]  & n8423;
  assign n8426 = ~n8424 & ~n8425;
  assign n8427 = ~n8407 & ~n8426;
  assign n8428 = n7982 & ~n7995;
  assign n8429 = ~n7994 & ~n7995;
  assign n8430 = ~n8428 & ~n8429;
  assign n8431 = n8407 & n8426;
  assign n8432 = ~n8427 & ~n8431;
  assign n8433 = ~n8430 & n8432;
  assign n8434 = ~n8427 & ~n8433;
  assign n8435 = ~n8021 & ~n8434;
  assign n8436 = n8021 & n8434;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = ~n8430 & ~n8433;
  assign n8439 = n8432 & ~n8433;
  assign n8440 = ~n8438 & ~n8439;
  assign n8441 = n8374 & ~n8386;
  assign n8442 = ~n8385 & ~n8386;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = n8358 & ~n8370;
  assign n8445 = ~n8369 & ~n8370;
  assign n8446 = ~n8444 & ~n8445;
  assign n8447 = n8062 & n8335;
  assign n8448 = ~n8336 & ~n8447;
  assign n8449 = ~n1235 & n5496;
  assign n8450 = ~n1472 & n4935;
  assign n8451 = ~n1364 & n5407;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = ~n8449 & n8452;
  assign n8454 = ~n4938 & n8453;
  assign n8455 = ~n4848 & n8453;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 =  a[20]  & ~n8456;
  assign n8458 = ~ a[20]  & n8456;
  assign n8459 = ~n8457 & ~n8458;
  assign n8460 = n8448 & ~n8459;
  assign n8461 = n8080 & n8333;
  assign n8462 = ~n8334 & ~n8461;
  assign n8463 = ~n1364 & n5496;
  assign n8464 = ~n1572 & n4935;
  assign n8465 = ~n1472 & n5407;
  assign n8466 = ~n8464 & ~n8465;
  assign n8467 = ~n8463 & n8466;
  assign n8468 = ~n4938 & n8467;
  assign n8469 = ~n5114 & n8467;
  assign n8470 = ~n8468 & ~n8469;
  assign n8471 =  a[20]  & ~n8470;
  assign n8472 = ~ a[20]  & n8470;
  assign n8473 = ~n8471 & ~n8472;
  assign n8474 = n8462 & ~n8473;
  assign n8475 = n8098 & n8331;
  assign n8476 = ~n8332 & ~n8475;
  assign n8477 = ~n1472 & n5496;
  assign n8478 = ~n1665 & n4935;
  assign n8479 = ~n1572 & n5407;
  assign n8480 = ~n8478 & ~n8479;
  assign n8481 = ~n8477 & n8480;
  assign n8482 = ~n4938 & n8481;
  assign n8483 = ~n5139 & n8481;
  assign n8484 = ~n8482 & ~n8483;
  assign n8485 =  a[20]  & ~n8484;
  assign n8486 = ~ a[20]  & n8484;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = n8476 & ~n8487;
  assign n8489 = n8116 & n8329;
  assign n8490 = ~n8330 & ~n8489;
  assign n8491 = ~n1572 & n5496;
  assign n8492 = ~n1779 & n4935;
  assign n8493 = ~n1665 & n5407;
  assign n8494 = ~n8492 & ~n8493;
  assign n8495 = ~n8491 & n8494;
  assign n8496 = ~n4938 & n8495;
  assign n8497 = ~n5561 & n8495;
  assign n8498 = ~n8496 & ~n8497;
  assign n8499 =  a[20]  & ~n8498;
  assign n8500 = ~ a[20]  & n8498;
  assign n8501 = ~n8499 & ~n8500;
  assign n8502 = n8490 & ~n8501;
  assign n8503 = n8134 & n8327;
  assign n8504 = ~n8328 & ~n8503;
  assign n8505 = ~n1665 & n5496;
  assign n8506 = ~n1877 & n4935;
  assign n8507 = ~n1779 & n5407;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = ~n8505 & n8508;
  assign n8510 = ~n4938 & n8509;
  assign n8511 = ~n5328 & n8509;
  assign n8512 = ~n8510 & ~n8511;
  assign n8513 =  a[20]  & ~n8512;
  assign n8514 = ~ a[20]  & n8512;
  assign n8515 = ~n8513 & ~n8514;
  assign n8516 = n8504 & ~n8515;
  assign n8517 = n8152 & n8325;
  assign n8518 = ~n8326 & ~n8517;
  assign n8519 = ~n1779 & n5496;
  assign n8520 = ~n1913 & n4935;
  assign n8521 = ~n1877 & n5407;
  assign n8522 = ~n8520 & ~n8521;
  assign n8523 = ~n8519 & n8522;
  assign n8524 = ~n4938 & n8523;
  assign n8525 = ~n5851 & n8523;
  assign n8526 = ~n8524 & ~n8525;
  assign n8527 =  a[20]  & ~n8526;
  assign n8528 = ~ a[20]  & n8526;
  assign n8529 = ~n8527 & ~n8528;
  assign n8530 = n8518 & ~n8529;
  assign n8531 = n8170 & n8323;
  assign n8532 = ~n8324 & ~n8531;
  assign n8533 = ~n1877 & n5496;
  assign n8534 = ~n1992 & n4935;
  assign n8535 = ~n1913 & n5407;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = ~n8533 & n8536;
  assign n8538 = ~n4938 & n8537;
  assign n8539 = ~n6007 & n8537;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 =  a[20]  & ~n8540;
  assign n8542 = ~ a[20]  & n8540;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = n8532 & ~n8543;
  assign n8545 = ~n1913 & n5496;
  assign n8546 = ~n2057 & n4935;
  assign n8547 = ~n1992 & n5407;
  assign n8548 = ~n8546 & ~n8547;
  assign n8549 = ~n8545 & n8548;
  assign n8550 = n4938 & n5834;
  assign n8551 = n8549 & ~n8550;
  assign n8552 =  a[20]  & ~n8551;
  assign n8553 = ~n8551 & ~n8552;
  assign n8554 =  a[20]  & ~n8552;
  assign n8555 = ~n8553 & ~n8554;
  assign n8556 = n8319 & ~n8321;
  assign n8557 = ~n8322 & ~n8556;
  assign n8558 = ~n8555 & n8557;
  assign n8559 = ~n8555 & ~n8558;
  assign n8560 = n8557 & ~n8558;
  assign n8561 = ~n8559 & ~n8560;
  assign n8562 = ~n1992 & n5496;
  assign n8563 = ~n2152 & n4935;
  assign n8564 = ~n2057 & n5407;
  assign n8565 = ~n8563 & ~n8564;
  assign n8566 = ~n8562 & n8565;
  assign n8567 = n4938 & n6143;
  assign n8568 = n8566 & ~n8567;
  assign n8569 =  a[20]  & ~n8568;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 =  a[20]  & ~n8569;
  assign n8572 = ~n8570 & ~n8571;
  assign n8573 = ~n8314 & ~n8318;
  assign n8574 = ~n8317 & ~n8318;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = ~n8572 & ~n8575;
  assign n8577 = ~n8572 & ~n8576;
  assign n8578 = ~n8575 & ~n8576;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = n8215 & n8312;
  assign n8581 = ~n8313 & ~n8580;
  assign n8582 = ~n2057 & n5496;
  assign n8583 = ~n2189 & n4935;
  assign n8584 = ~n2152 & n5407;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = ~n8582 & n8585;
  assign n8587 = ~n4938 & n8586;
  assign n8588 = ~n6479 & n8586;
  assign n8589 = ~n8587 & ~n8588;
  assign n8590 =  a[20]  & ~n8589;
  assign n8591 = ~ a[20]  & n8589;
  assign n8592 = ~n8590 & ~n8591;
  assign n8593 = n8581 & ~n8592;
  assign n8594 = n8308 & ~n8310;
  assign n8595 = ~n8311 & ~n8594;
  assign n8596 = ~n2152 & n5496;
  assign n8597 = ~n2291 & n4935;
  assign n8598 = ~n2189 & n5407;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = ~n8596 & n8599;
  assign n8601 = ~n4938 & n8600;
  assign n8602 = ~n6492 & n8600;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 =  a[20]  & ~n8603;
  assign n8605 = ~ a[20]  & n8603;
  assign n8606 = ~n8604 & ~n8605;
  assign n8607 = n8595 & ~n8606;
  assign n8608 = n8247 & n8306;
  assign n8609 = ~n8307 & ~n8608;
  assign n8610 = ~n2189 & n5496;
  assign n8611 = ~n2388 & n4935;
  assign n8612 = ~n2291 & n5407;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = ~n8610 & n8613;
  assign n8615 = ~n4938 & n8614;
  assign n8616 = ~n6122 & n8614;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 =  a[20]  & ~n8617;
  assign n8619 = ~ a[20]  & n8617;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = n8609 & ~n8620;
  assign n8622 = ~n2291 & n5496;
  assign n8623 = ~n2464 & n4935;
  assign n8624 = ~n2388 & n5407;
  assign n8625 = ~n8623 & ~n8624;
  assign n8626 = ~n8622 & n8625;
  assign n8627 = n4938 & n6541;
  assign n8628 = n8626 & ~n8627;
  assign n8629 =  a[20]  & ~n8628;
  assign n8630 = ~n8628 & ~n8629;
  assign n8631 =  a[20]  & ~n8629;
  assign n8632 = ~n8630 & ~n8631;
  assign n8633 = n8302 & ~n8304;
  assign n8634 = ~n8305 & ~n8633;
  assign n8635 = ~n8632 & n8634;
  assign n8636 = ~n8632 & ~n8635;
  assign n8637 = n8634 & ~n8635;
  assign n8638 = ~n8636 & ~n8637;
  assign n8639 = ~n8289 & ~n8301;
  assign n8640 = ~n8300 & ~n8301;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = ~n2388 & n5496;
  assign n8643 = ~n2533 & n4935;
  assign n8644 = ~n2464 & n5407;
  assign n8645 = ~n8643 & ~n8644;
  assign n8646 = ~n8642 & n8645;
  assign n8647 = ~n4938 & n8646;
  assign n8648 = ~n6591 & n8646;
  assign n8649 = ~n8647 & ~n8648;
  assign n8650 =  a[20]  & ~n8649;
  assign n8651 = ~ a[20]  & n8649;
  assign n8652 = ~n8650 & ~n8651;
  assign n8653 = ~n8641 & ~n8652;
  assign n8654 = ~n2464 & n5496;
  assign n8655 = ~n2571 & n4935;
  assign n8656 = ~n2533 & n5407;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = ~n8654 & n8657;
  assign n8659 = n4938 & n6646;
  assign n8660 = n8658 & ~n8659;
  assign n8661 =  a[20]  & ~n8660;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 =  a[20]  & ~n8661;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = ~n8273 & n8284;
  assign n8666 = ~n8285 & ~n8665;
  assign n8667 = ~n8664 & n8666;
  assign n8668 = ~n8664 & ~n8667;
  assign n8669 = n8666 & ~n8667;
  assign n8670 = ~n8668 & ~n8669;
  assign n8671 = n8270 & ~n8272;
  assign n8672 = ~n8273 & ~n8671;
  assign n8673 = ~n2533 & n5496;
  assign n8674 = ~n2674 & n4935;
  assign n8675 = ~n2571 & n5407;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = ~n8673 & n8676;
  assign n8678 = ~n4938 & n8677;
  assign n8679 = ~n6695 & n8677;
  assign n8680 = ~n8678 & ~n8679;
  assign n8681 =  a[20]  & ~n8680;
  assign n8682 = ~ a[20]  & n8680;
  assign n8683 = ~n8681 & ~n8682;
  assign n8684 = n8672 & ~n8683;
  assign n8685 = ~n2829 & n5407;
  assign n8686 = ~n2736 & n5496;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = n4938 & ~n7469;
  assign n8689 = n8687 & ~n8688;
  assign n8690 =  a[20]  & ~n8689;
  assign n8691 =  a[20]  & ~n8690;
  assign n8692 = ~n8689 & ~n8690;
  assign n8693 = ~n8691 & ~n8692;
  assign n8694 = ~n2829 & ~n4933;
  assign n8695 =  a[20]  & ~n8694;
  assign n8696 = ~n8693 & n8695;
  assign n8697 = ~n2674 & n5496;
  assign n8698 = ~n2829 & n4935;
  assign n8699 = ~n2736 & n5407;
  assign n8700 = ~n8698 & ~n8699;
  assign n8701 = ~n8697 & n8700;
  assign n8702 = ~n4938 & n8701;
  assign n8703 = ~n6798 & n8701;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 =  a[20]  & ~n8704;
  assign n8706 = ~ a[20]  & n8704;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = n8696 & ~n8707;
  assign n8709 = n8271 & n8708;
  assign n8710 = n8708 & ~n8709;
  assign n8711 = n8271 & ~n8709;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = ~n2571 & n5496;
  assign n8714 = ~n2736 & n4935;
  assign n8715 = ~n2674 & n5407;
  assign n8716 = ~n8714 & ~n8715;
  assign n8717 = ~n8713 & n8716;
  assign n8718 = n4938 & n6806;
  assign n8719 = n8717 & ~n8718;
  assign n8720 =  a[20]  & ~n8719;
  assign n8721 =  a[20]  & ~n8720;
  assign n8722 = ~n8719 & ~n8720;
  assign n8723 = ~n8721 & ~n8722;
  assign n8724 = ~n8712 & ~n8723;
  assign n8725 = ~n8709 & ~n8724;
  assign n8726 = ~n8672 & n8683;
  assign n8727 = ~n8684 & ~n8726;
  assign n8728 = ~n8725 & n8727;
  assign n8729 = ~n8684 & ~n8728;
  assign n8730 = ~n8670 & ~n8729;
  assign n8731 = ~n8667 & ~n8730;
  assign n8732 = n8641 & n8652;
  assign n8733 = ~n8653 & ~n8732;
  assign n8734 = ~n8731 & n8733;
  assign n8735 = ~n8653 & ~n8734;
  assign n8736 = ~n8638 & ~n8735;
  assign n8737 = ~n8635 & ~n8736;
  assign n8738 = n8609 & ~n8621;
  assign n8739 = ~n8620 & ~n8621;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~n8737 & ~n8740;
  assign n8742 = ~n8621 & ~n8741;
  assign n8743 = n8595 & ~n8607;
  assign n8744 = ~n8606 & ~n8607;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = ~n8742 & ~n8745;
  assign n8747 = ~n8607 & ~n8746;
  assign n8748 = ~n8581 & n8592;
  assign n8749 = ~n8593 & ~n8748;
  assign n8750 = ~n8747 & n8749;
  assign n8751 = ~n8593 & ~n8750;
  assign n8752 = ~n8579 & ~n8751;
  assign n8753 = ~n8576 & ~n8752;
  assign n8754 = ~n8561 & ~n8753;
  assign n8755 = ~n8558 & ~n8754;
  assign n8756 = n8532 & ~n8544;
  assign n8757 = ~n8543 & ~n8544;
  assign n8758 = ~n8756 & ~n8757;
  assign n8759 = ~n8755 & ~n8758;
  assign n8760 = ~n8544 & ~n8759;
  assign n8761 = n8518 & ~n8530;
  assign n8762 = ~n8529 & ~n8530;
  assign n8763 = ~n8761 & ~n8762;
  assign n8764 = ~n8760 & ~n8763;
  assign n8765 = ~n8530 & ~n8764;
  assign n8766 = n8504 & ~n8516;
  assign n8767 = ~n8515 & ~n8516;
  assign n8768 = ~n8766 & ~n8767;
  assign n8769 = ~n8765 & ~n8768;
  assign n8770 = ~n8516 & ~n8769;
  assign n8771 = n8490 & ~n8502;
  assign n8772 = ~n8501 & ~n8502;
  assign n8773 = ~n8771 & ~n8772;
  assign n8774 = ~n8770 & ~n8773;
  assign n8775 = ~n8502 & ~n8774;
  assign n8776 = n8476 & ~n8488;
  assign n8777 = ~n8487 & ~n8488;
  assign n8778 = ~n8776 & ~n8777;
  assign n8779 = ~n8775 & ~n8778;
  assign n8780 = ~n8488 & ~n8779;
  assign n8781 = n8462 & ~n8474;
  assign n8782 = ~n8473 & ~n8474;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = ~n8780 & ~n8783;
  assign n8785 = ~n8474 & ~n8784;
  assign n8786 = n8448 & ~n8460;
  assign n8787 = ~n8459 & ~n8460;
  assign n8788 = ~n8786 & ~n8787;
  assign n8789 = ~n8785 & ~n8788;
  assign n8790 = ~n8460 & ~n8789;
  assign n8791 = n8351 & ~n8353;
  assign n8792 = ~n8354 & ~n8791;
  assign n8793 = ~n8790 & n8792;
  assign n8794 = ~n867 & n6233;
  assign n8795 = ~n1060 & n5663;
  assign n8796 = ~n958 & n5939;
  assign n8797 = ~n8795 & ~n8796;
  assign n8798 = ~n8794 & n8797;
  assign n8799 = n4204 & n5666;
  assign n8800 = n8798 & ~n8799;
  assign n8801 =  a[17]  & ~n8800;
  assign n8802 = ~n8800 & ~n8801;
  assign n8803 =  a[17]  & ~n8801;
  assign n8804 = ~n8802 & ~n8803;
  assign n8805 = n8790 & ~n8792;
  assign n8806 = ~n8793 & ~n8805;
  assign n8807 = ~n8804 & n8806;
  assign n8808 = ~n8793 & ~n8807;
  assign n8809 = ~n8446 & ~n8808;
  assign n8810 = n8446 & n8808;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = ~n3012 & n7101;
  assign n8813 = ~n587 & n6402;
  assign n8814 = ~n392 & n6951;
  assign n8815 = ~n8813 & ~n8814;
  assign n8816 = ~n8812 & n8815;
  assign n8817 = n3018 & n6397;
  assign n8818 = n8816 & ~n8817;
  assign n8819 =  a[14]  & ~n8818;
  assign n8820 =  a[14]  & ~n8819;
  assign n8821 = ~n8818 & ~n8819;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = n8811 & ~n8822;
  assign n8824 = ~n8809 & ~n8823;
  assign n8825 = ~n8443 & ~n8824;
  assign n8826 = n8443 & n8824;
  assign n8827 = ~n8825 & ~n8826;
  assign n8828 = ~n3805 & n7983;
  assign n8829 = ~n3605 & n7291;
  assign n8830 = ~n3456 & n7632;
  assign n8831 = ~n8829 & ~n8830;
  assign n8832 = ~n8828 & n8831;
  assign n8833 = n3818 & n7294;
  assign n8834 = n8832 & ~n8833;
  assign n8835 =  a[11]  & ~n8834;
  assign n8836 =  a[11]  & ~n8835;
  assign n8837 = ~n8834 & ~n8835;
  assign n8838 = ~n8836 & ~n8837;
  assign n8839 = n8827 & ~n8838;
  assign n8840 = ~n8825 & ~n8839;
  assign n8841 = ~n3964 & n7983;
  assign n8842 = ~n3456 & n7291;
  assign n8843 = ~n3805 & n7632;
  assign n8844 = ~n8842 & ~n8843;
  assign n8845 = ~n8841 & n8844;
  assign n8846 = ~n7294 & n8845;
  assign n8847 = ~n4558 & n8845;
  assign n8848 = ~n8846 & ~n8847;
  assign n8849 =  a[11]  & ~n8848;
  assign n8850 = ~ a[11]  & n8848;
  assign n8851 = ~n8849 & ~n8850;
  assign n8852 = ~n8840 & ~n8851;
  assign n8853 = n8840 & n8851;
  assign n8854 = ~n8852 & ~n8853;
  assign n8855 = n8387 & ~n8389;
  assign n8856 = ~n8390 & ~n8855;
  assign n8857 = n8854 & n8856;
  assign n8858 = ~n8852 & ~n8857;
  assign n8859 = ~n3877 & n8418;
  assign n8860 = ~n8410 & n8416;
  assign n8861 = ~n4515 & n8860;
  assign n8862 = ~n8859 & ~n8861;
  assign n8863 = ~n8421 & n8862;
  assign n8864 = ~n4609 & n8862;
  assign n8865 = ~n8863 & ~n8864;
  assign n8866 =  a[8]  & ~n8865;
  assign n8867 = ~ a[8]  & n8865;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~n8858 & ~n8868;
  assign n8870 = n8394 & ~n8406;
  assign n8871 = ~n8405 & ~n8406;
  assign n8872 = ~n8870 & ~n8871;
  assign n8873 = n8858 & n8868;
  assign n8874 = ~n8869 & ~n8873;
  assign n8875 = ~n8872 & n8874;
  assign n8876 = ~n8869 & ~n8875;
  assign n8877 = ~n8440 & ~n8876;
  assign n8878 = n8440 & n8876;
  assign n8879 = ~n8877 & ~n8878;
  assign n8880 = n8827 & ~n8839;
  assign n8881 = ~n8838 & ~n8839;
  assign n8882 = ~n8880 & ~n8881;
  assign n8883 = n8811 & ~n8823;
  assign n8884 = ~n8822 & ~n8823;
  assign n8885 = ~n8883 & ~n8884;
  assign n8886 = ~n958 & n6233;
  assign n8887 = ~n1178 & n5663;
  assign n8888 = ~n1060 & n5939;
  assign n8889 = ~n8887 & ~n8888;
  assign n8890 = ~n8886 & n8889;
  assign n8891 = n4633 & n5666;
  assign n8892 = n8890 & ~n8891;
  assign n8893 =  a[17]  & ~n8892;
  assign n8894 = ~n8892 & ~n8893;
  assign n8895 =  a[17]  & ~n8893;
  assign n8896 = ~n8894 & ~n8895;
  assign n8897 = ~n8785 & ~n8789;
  assign n8898 = ~n8788 & ~n8789;
  assign n8899 = ~n8897 & ~n8898;
  assign n8900 = ~n8896 & ~n8899;
  assign n8901 = ~n8896 & ~n8900;
  assign n8902 = ~n8899 & ~n8900;
  assign n8903 = ~n8901 & ~n8902;
  assign n8904 = ~n1060 & n6233;
  assign n8905 = ~n1235 & n5663;
  assign n8906 = ~n1178 & n5939;
  assign n8907 = ~n8905 & ~n8906;
  assign n8908 = ~n8904 & n8907;
  assign n8909 = n4429 & n5666;
  assign n8910 = n8908 & ~n8909;
  assign n8911 =  a[17]  & ~n8910;
  assign n8912 = ~n8910 & ~n8911;
  assign n8913 =  a[17]  & ~n8911;
  assign n8914 = ~n8912 & ~n8913;
  assign n8915 = ~n8780 & ~n8784;
  assign n8916 = ~n8783 & ~n8784;
  assign n8917 = ~n8915 & ~n8916;
  assign n8918 = ~n8914 & ~n8917;
  assign n8919 = ~n8914 & ~n8918;
  assign n8920 = ~n8917 & ~n8918;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = ~n1178 & n6233;
  assign n8923 = ~n1364 & n5663;
  assign n8924 = ~n1235 & n5939;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = ~n8922 & n8925;
  assign n8927 = n4861 & n5666;
  assign n8928 = n8926 & ~n8927;
  assign n8929 =  a[17]  & ~n8928;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 =  a[17]  & ~n8929;
  assign n8932 = ~n8930 & ~n8931;
  assign n8933 = ~n8775 & ~n8779;
  assign n8934 = ~n8778 & ~n8779;
  assign n8935 = ~n8933 & ~n8934;
  assign n8936 = ~n8932 & ~n8935;
  assign n8937 = ~n8932 & ~n8936;
  assign n8938 = ~n8935 & ~n8936;
  assign n8939 = ~n8937 & ~n8938;
  assign n8940 = ~n1235 & n6233;
  assign n8941 = ~n1472 & n5663;
  assign n8942 = ~n1364 & n5939;
  assign n8943 = ~n8941 & ~n8942;
  assign n8944 = ~n8940 & n8943;
  assign n8945 = n4848 & n5666;
  assign n8946 = n8944 & ~n8945;
  assign n8947 =  a[17]  & ~n8946;
  assign n8948 = ~n8946 & ~n8947;
  assign n8949 =  a[17]  & ~n8947;
  assign n8950 = ~n8948 & ~n8949;
  assign n8951 = ~n8770 & ~n8774;
  assign n8952 = ~n8773 & ~n8774;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = ~n8950 & ~n8953;
  assign n8955 = ~n8950 & ~n8954;
  assign n8956 = ~n8953 & ~n8954;
  assign n8957 = ~n8955 & ~n8956;
  assign n8958 = ~n1364 & n6233;
  assign n8959 = ~n1572 & n5663;
  assign n8960 = ~n1472 & n5939;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = ~n8958 & n8961;
  assign n8963 = n5114 & n5666;
  assign n8964 = n8962 & ~n8963;
  assign n8965 =  a[17]  & ~n8964;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 =  a[17]  & ~n8965;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = ~n8765 & ~n8769;
  assign n8970 = ~n8768 & ~n8769;
  assign n8971 = ~n8969 & ~n8970;
  assign n8972 = ~n8968 & ~n8971;
  assign n8973 = ~n8968 & ~n8972;
  assign n8974 = ~n8971 & ~n8972;
  assign n8975 = ~n8973 & ~n8974;
  assign n8976 = ~n1472 & n6233;
  assign n8977 = ~n1665 & n5663;
  assign n8978 = ~n1572 & n5939;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = ~n8976 & n8979;
  assign n8981 = n5139 & n5666;
  assign n8982 = n8980 & ~n8981;
  assign n8983 =  a[17]  & ~n8982;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 =  a[17]  & ~n8983;
  assign n8986 = ~n8984 & ~n8985;
  assign n8987 = ~n8760 & ~n8764;
  assign n8988 = ~n8763 & ~n8764;
  assign n8989 = ~n8987 & ~n8988;
  assign n8990 = ~n8986 & ~n8989;
  assign n8991 = ~n8986 & ~n8990;
  assign n8992 = ~n8989 & ~n8990;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = ~n1572 & n6233;
  assign n8995 = ~n1779 & n5663;
  assign n8996 = ~n1665 & n5939;
  assign n8997 = ~n8995 & ~n8996;
  assign n8998 = ~n8994 & n8997;
  assign n8999 = n5561 & n5666;
  assign n9000 = n8998 & ~n8999;
  assign n9001 =  a[17]  & ~n9000;
  assign n9002 = ~n9000 & ~n9001;
  assign n9003 =  a[17]  & ~n9001;
  assign n9004 = ~n9002 & ~n9003;
  assign n9005 = ~n8755 & ~n8759;
  assign n9006 = ~n8758 & ~n8759;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = ~n9004 & ~n9007;
  assign n9009 = ~n9004 & ~n9008;
  assign n9010 = ~n9007 & ~n9008;
  assign n9011 = ~n9009 & ~n9010;
  assign n9012 = n8561 & n8753;
  assign n9013 = ~n8754 & ~n9012;
  assign n9014 = ~n1665 & n6233;
  assign n9015 = ~n1877 & n5663;
  assign n9016 = ~n1779 & n5939;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = ~n9014 & n9017;
  assign n9019 = ~n5666 & n9018;
  assign n9020 = ~n5328 & n9018;
  assign n9021 = ~n9019 & ~n9020;
  assign n9022 =  a[17]  & ~n9021;
  assign n9023 = ~ a[17]  & n9021;
  assign n9024 = ~n9022 & ~n9023;
  assign n9025 = n9013 & ~n9024;
  assign n9026 = n8579 & n8751;
  assign n9027 = ~n8752 & ~n9026;
  assign n9028 = ~n1779 & n6233;
  assign n9029 = ~n1913 & n5663;
  assign n9030 = ~n1877 & n5939;
  assign n9031 = ~n9029 & ~n9030;
  assign n9032 = ~n9028 & n9031;
  assign n9033 = ~n5666 & n9032;
  assign n9034 = ~n5851 & n9032;
  assign n9035 = ~n9033 & ~n9034;
  assign n9036 =  a[17]  & ~n9035;
  assign n9037 = ~ a[17]  & n9035;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = n9027 & ~n9038;
  assign n9040 = ~n1877 & n6233;
  assign n9041 = ~n1992 & n5663;
  assign n9042 = ~n1913 & n5939;
  assign n9043 = ~n9041 & ~n9042;
  assign n9044 = ~n9040 & n9043;
  assign n9045 = n5666 & n6007;
  assign n9046 = n9044 & ~n9045;
  assign n9047 =  a[17]  & ~n9046;
  assign n9048 = ~n9046 & ~n9047;
  assign n9049 =  a[17]  & ~n9047;
  assign n9050 = ~n9048 & ~n9049;
  assign n9051 = n8747 & ~n8749;
  assign n9052 = ~n8750 & ~n9051;
  assign n9053 = ~n9050 & n9052;
  assign n9054 = ~n9050 & ~n9053;
  assign n9055 = n9052 & ~n9053;
  assign n9056 = ~n9054 & ~n9055;
  assign n9057 = ~n1913 & n6233;
  assign n9058 = ~n2057 & n5663;
  assign n9059 = ~n1992 & n5939;
  assign n9060 = ~n9058 & ~n9059;
  assign n9061 = ~n9057 & n9060;
  assign n9062 = n5666 & n5834;
  assign n9063 = n9061 & ~n9062;
  assign n9064 =  a[17]  & ~n9063;
  assign n9065 = ~n9063 & ~n9064;
  assign n9066 =  a[17]  & ~n9064;
  assign n9067 = ~n9065 & ~n9066;
  assign n9068 = ~n8742 & ~n8746;
  assign n9069 = ~n8745 & ~n8746;
  assign n9070 = ~n9068 & ~n9069;
  assign n9071 = ~n9067 & ~n9070;
  assign n9072 = ~n9067 & ~n9071;
  assign n9073 = ~n9070 & ~n9071;
  assign n9074 = ~n9072 & ~n9073;
  assign n9075 = ~n1992 & n6233;
  assign n9076 = ~n2152 & n5663;
  assign n9077 = ~n2057 & n5939;
  assign n9078 = ~n9076 & ~n9077;
  assign n9079 = ~n9075 & n9078;
  assign n9080 = n5666 & n6143;
  assign n9081 = n9079 & ~n9080;
  assign n9082 =  a[17]  & ~n9081;
  assign n9083 = ~n9081 & ~n9082;
  assign n9084 =  a[17]  & ~n9082;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = ~n8737 & ~n8741;
  assign n9087 = ~n8740 & ~n8741;
  assign n9088 = ~n9086 & ~n9087;
  assign n9089 = ~n9085 & ~n9088;
  assign n9090 = ~n9085 & ~n9089;
  assign n9091 = ~n9088 & ~n9089;
  assign n9092 = ~n9090 & ~n9091;
  assign n9093 = n8638 & n8735;
  assign n9094 = ~n8736 & ~n9093;
  assign n9095 = ~n2057 & n6233;
  assign n9096 = ~n2189 & n5663;
  assign n9097 = ~n2152 & n5939;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = ~n9095 & n9098;
  assign n9100 = ~n5666 & n9099;
  assign n9101 = ~n6479 & n9099;
  assign n9102 = ~n9100 & ~n9101;
  assign n9103 =  a[17]  & ~n9102;
  assign n9104 = ~ a[17]  & n9102;
  assign n9105 = ~n9103 & ~n9104;
  assign n9106 = n9094 & ~n9105;
  assign n9107 = n8731 & ~n8733;
  assign n9108 = ~n8734 & ~n9107;
  assign n9109 = ~n2152 & n6233;
  assign n9110 = ~n2291 & n5663;
  assign n9111 = ~n2189 & n5939;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = ~n9109 & n9112;
  assign n9114 = ~n5666 & n9113;
  assign n9115 = ~n6492 & n9113;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 =  a[17]  & ~n9116;
  assign n9118 = ~ a[17]  & n9116;
  assign n9119 = ~n9117 & ~n9118;
  assign n9120 = n9108 & ~n9119;
  assign n9121 = n8670 & n8729;
  assign n9122 = ~n8730 & ~n9121;
  assign n9123 = ~n2189 & n6233;
  assign n9124 = ~n2388 & n5663;
  assign n9125 = ~n2291 & n5939;
  assign n9126 = ~n9124 & ~n9125;
  assign n9127 = ~n9123 & n9126;
  assign n9128 = ~n5666 & n9127;
  assign n9129 = ~n6122 & n9127;
  assign n9130 = ~n9128 & ~n9129;
  assign n9131 =  a[17]  & ~n9130;
  assign n9132 = ~ a[17]  & n9130;
  assign n9133 = ~n9131 & ~n9132;
  assign n9134 = n9122 & ~n9133;
  assign n9135 = ~n2291 & n6233;
  assign n9136 = ~n2464 & n5663;
  assign n9137 = ~n2388 & n5939;
  assign n9138 = ~n9136 & ~n9137;
  assign n9139 = ~n9135 & n9138;
  assign n9140 = n5666 & n6541;
  assign n9141 = n9139 & ~n9140;
  assign n9142 =  a[17]  & ~n9141;
  assign n9143 = ~n9141 & ~n9142;
  assign n9144 =  a[17]  & ~n9142;
  assign n9145 = ~n9143 & ~n9144;
  assign n9146 = n8725 & ~n8727;
  assign n9147 = ~n8728 & ~n9146;
  assign n9148 = ~n9145 & n9147;
  assign n9149 = ~n9145 & ~n9148;
  assign n9150 = n9147 & ~n9148;
  assign n9151 = ~n9149 & ~n9150;
  assign n9152 = ~n8712 & ~n8724;
  assign n9153 = ~n8723 & ~n8724;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = ~n2388 & n6233;
  assign n9156 = ~n2533 & n5663;
  assign n9157 = ~n2464 & n5939;
  assign n9158 = ~n9156 & ~n9157;
  assign n9159 = ~n9155 & n9158;
  assign n9160 = ~n5666 & n9159;
  assign n9161 = ~n6591 & n9159;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 =  a[17]  & ~n9162;
  assign n9164 = ~ a[17]  & n9162;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = ~n9154 & ~n9165;
  assign n9167 = ~n2464 & n6233;
  assign n9168 = ~n2571 & n5663;
  assign n9169 = ~n2533 & n5939;
  assign n9170 = ~n9168 & ~n9169;
  assign n9171 = ~n9167 & n9170;
  assign n9172 = n5666 & n6646;
  assign n9173 = n9171 & ~n9172;
  assign n9174 =  a[17]  & ~n9173;
  assign n9175 = ~n9173 & ~n9174;
  assign n9176 =  a[17]  & ~n9174;
  assign n9177 = ~n9175 & ~n9176;
  assign n9178 = ~n8696 & n8707;
  assign n9179 = ~n8708 & ~n9178;
  assign n9180 = ~n9177 & n9179;
  assign n9181 = ~n9177 & ~n9180;
  assign n9182 = n9179 & ~n9180;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = n8693 & ~n8695;
  assign n9185 = ~n8696 & ~n9184;
  assign n9186 = ~n2533 & n6233;
  assign n9187 = ~n2674 & n5663;
  assign n9188 = ~n2571 & n5939;
  assign n9189 = ~n9187 & ~n9188;
  assign n9190 = ~n9186 & n9189;
  assign n9191 = ~n5666 & n9190;
  assign n9192 = ~n6695 & n9190;
  assign n9193 = ~n9191 & ~n9192;
  assign n9194 =  a[17]  & ~n9193;
  assign n9195 = ~ a[17]  & n9193;
  assign n9196 = ~n9194 & ~n9195;
  assign n9197 = n9185 & ~n9196;
  assign n9198 = ~n2829 & n5939;
  assign n9199 = ~n2736 & n6233;
  assign n9200 = ~n9198 & ~n9199;
  assign n9201 = n5666 & ~n7469;
  assign n9202 = n9200 & ~n9201;
  assign n9203 =  a[17]  & ~n9202;
  assign n9204 =  a[17]  & ~n9203;
  assign n9205 = ~n9202 & ~n9203;
  assign n9206 = ~n9204 & ~n9205;
  assign n9207 = ~n2829 & ~n5658;
  assign n9208 =  a[17]  & ~n9207;
  assign n9209 = ~n9206 & n9208;
  assign n9210 = ~n2674 & n6233;
  assign n9211 = ~n2829 & n5663;
  assign n9212 = ~n2736 & n5939;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~n9210 & n9213;
  assign n9215 = ~n5666 & n9214;
  assign n9216 = ~n6798 & n9214;
  assign n9217 = ~n9215 & ~n9216;
  assign n9218 =  a[17]  & ~n9217;
  assign n9219 = ~ a[17]  & n9217;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = n9209 & ~n9220;
  assign n9222 = n8694 & n9221;
  assign n9223 = n9221 & ~n9222;
  assign n9224 = n8694 & ~n9222;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = ~n2571 & n6233;
  assign n9227 = ~n2736 & n5663;
  assign n9228 = ~n2674 & n5939;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = ~n9226 & n9229;
  assign n9231 = n5666 & n6806;
  assign n9232 = n9230 & ~n9231;
  assign n9233 =  a[17]  & ~n9232;
  assign n9234 =  a[17]  & ~n9233;
  assign n9235 = ~n9232 & ~n9233;
  assign n9236 = ~n9234 & ~n9235;
  assign n9237 = ~n9225 & ~n9236;
  assign n9238 = ~n9222 & ~n9237;
  assign n9239 = ~n9185 & n9196;
  assign n9240 = ~n9197 & ~n9239;
  assign n9241 = ~n9238 & n9240;
  assign n9242 = ~n9197 & ~n9241;
  assign n9243 = ~n9183 & ~n9242;
  assign n9244 = ~n9180 & ~n9243;
  assign n9245 = n9154 & n9165;
  assign n9246 = ~n9166 & ~n9245;
  assign n9247 = ~n9244 & n9246;
  assign n9248 = ~n9166 & ~n9247;
  assign n9249 = ~n9151 & ~n9248;
  assign n9250 = ~n9148 & ~n9249;
  assign n9251 = n9122 & ~n9134;
  assign n9252 = ~n9133 & ~n9134;
  assign n9253 = ~n9251 & ~n9252;
  assign n9254 = ~n9250 & ~n9253;
  assign n9255 = ~n9134 & ~n9254;
  assign n9256 = n9108 & ~n9120;
  assign n9257 = ~n9119 & ~n9120;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = ~n9255 & ~n9258;
  assign n9260 = ~n9120 & ~n9259;
  assign n9261 = ~n9094 & n9105;
  assign n9262 = ~n9106 & ~n9261;
  assign n9263 = ~n9260 & n9262;
  assign n9264 = ~n9106 & ~n9263;
  assign n9265 = ~n9092 & ~n9264;
  assign n9266 = ~n9089 & ~n9265;
  assign n9267 = ~n9074 & ~n9266;
  assign n9268 = ~n9071 & ~n9267;
  assign n9269 = ~n9056 & ~n9268;
  assign n9270 = ~n9053 & ~n9269;
  assign n9271 = n9027 & ~n9039;
  assign n9272 = ~n9038 & ~n9039;
  assign n9273 = ~n9271 & ~n9272;
  assign n9274 = ~n9270 & ~n9273;
  assign n9275 = ~n9039 & ~n9274;
  assign n9276 = ~n9013 & n9024;
  assign n9277 = ~n9025 & ~n9276;
  assign n9278 = ~n9275 & n9277;
  assign n9279 = ~n9025 & ~n9278;
  assign n9280 = ~n9011 & ~n9279;
  assign n9281 = ~n9008 & ~n9280;
  assign n9282 = ~n8993 & ~n9281;
  assign n9283 = ~n8990 & ~n9282;
  assign n9284 = ~n8975 & ~n9283;
  assign n9285 = ~n8972 & ~n9284;
  assign n9286 = ~n8957 & ~n9285;
  assign n9287 = ~n8954 & ~n9286;
  assign n9288 = ~n8939 & ~n9287;
  assign n9289 = ~n8936 & ~n9288;
  assign n9290 = ~n8921 & ~n9289;
  assign n9291 = ~n8918 & ~n9290;
  assign n9292 = ~n8903 & ~n9291;
  assign n9293 = ~n8900 & ~n9292;
  assign n9294 = n8804 & ~n8806;
  assign n9295 = ~n8807 & ~n9294;
  assign n9296 = ~n9293 & n9295;
  assign n9297 = ~n392 & n7101;
  assign n9298 = ~n710 & n6402;
  assign n9299 = ~n587 & n6951;
  assign n9300 = ~n9298 & ~n9299;
  assign n9301 = ~n9297 & n9300;
  assign n9302 = n3347 & n6397;
  assign n9303 = n9301 & ~n9302;
  assign n9304 =  a[14]  & ~n9303;
  assign n9305 = ~n9303 & ~n9304;
  assign n9306 =  a[14]  & ~n9304;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = n9293 & ~n9295;
  assign n9309 = ~n9296 & ~n9308;
  assign n9310 = ~n9307 & n9309;
  assign n9311 = ~n9296 & ~n9310;
  assign n9312 = ~n8885 & ~n9311;
  assign n9313 = n8885 & n9311;
  assign n9314 = ~n9312 & ~n9313;
  assign n9315 = ~n3456 & n7983;
  assign n9316 = ~n3539 & n7291;
  assign n9317 = ~n3605 & n7632;
  assign n9318 = ~n9316 & ~n9317;
  assign n9319 = ~n9315 & n9318;
  assign n9320 = n3627 & n7294;
  assign n9321 = n9319 & ~n9320;
  assign n9322 =  a[11]  & ~n9321;
  assign n9323 =  a[11]  & ~n9322;
  assign n9324 = ~n9321 & ~n9322;
  assign n9325 = ~n9323 & ~n9324;
  assign n9326 = n9314 & ~n9325;
  assign n9327 = ~n9312 & ~n9326;
  assign n9328 = ~n8882 & ~n9327;
  assign n9329 = n8882 & n9327;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = n8413 & ~n8416;
  assign n9332 = ~n3877 & n9331;
  assign n9333 = ~n3964 & n8418;
  assign n9334 = ~n4045 & n8860;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = ~n9332 & n9335;
  assign n9337 = n4067 & n8421;
  assign n9338 = n9336 & ~n9337;
  assign n9339 =  a[8]  & ~n9338;
  assign n9340 =  a[8]  & ~n9339;
  assign n9341 = ~n9338 & ~n9339;
  assign n9342 = ~n9340 & ~n9341;
  assign n9343 = n9330 & ~n9342;
  assign n9344 = ~n9328 & ~n9343;
  assign n9345 = ~n4515 & n9331;
  assign n9346 = ~n4045 & n8418;
  assign n9347 = ~n3877 & n8860;
  assign n9348 = ~n9346 & ~n9347;
  assign n9349 = ~n9345 & n9348;
  assign n9350 = ~n8421 & n9349;
  assign n9351 = ~n4715 & n9349;
  assign n9352 = ~n9350 & ~n9351;
  assign n9353 =  a[8]  & ~n9352;
  assign n9354 = ~ a[8]  & n9352;
  assign n9355 = ~n9353 & ~n9354;
  assign n9356 = ~n9344 & ~n9355;
  assign n9357 = ~n9344 & ~n9356;
  assign n9358 = ~n9355 & ~n9356;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = ~n8854 & ~n8856;
  assign n9361 = ~n8857 & ~n9360;
  assign n9362 = ~n9359 & n9361;
  assign n9363 = ~n9356 & ~n9362;
  assign n9364 = n8872 & ~n8874;
  assign n9365 = ~n8875 & ~n9364;
  assign n9366 = ~n9363 & n9365;
  assign n9367 = n9314 & ~n9326;
  assign n9368 = ~n9325 & ~n9326;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = n8903 & n9291;
  assign n9371 = ~n9292 & ~n9370;
  assign n9372 = ~n587 & n7101;
  assign n9373 = ~n867 & n6402;
  assign n9374 = ~n710 & n6951;
  assign n9375 = ~n9373 & ~n9374;
  assign n9376 = ~n9372 & n9375;
  assign n9377 = ~n6397 & n9376;
  assign n9378 = ~n3331 & n9376;
  assign n9379 = ~n9377 & ~n9378;
  assign n9380 =  a[14]  & ~n9379;
  assign n9381 = ~ a[14]  & n9379;
  assign n9382 = ~n9380 & ~n9381;
  assign n9383 = n9371 & ~n9382;
  assign n9384 = n8921 & n9289;
  assign n9385 = ~n9290 & ~n9384;
  assign n9386 = ~n710 & n7101;
  assign n9387 = ~n958 & n6402;
  assign n9388 = ~n867 & n6951;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = ~n9386 & n9389;
  assign n9391 = ~n6397 & n9390;
  assign n9392 = ~n4179 & n9390;
  assign n9393 = ~n9391 & ~n9392;
  assign n9394 =  a[14]  & ~n9393;
  assign n9395 = ~ a[14]  & n9393;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = n9385 & ~n9396;
  assign n9398 = n8939 & n9287;
  assign n9399 = ~n9288 & ~n9398;
  assign n9400 = ~n867 & n7101;
  assign n9401 = ~n1060 & n6402;
  assign n9402 = ~n958 & n6951;
  assign n9403 = ~n9401 & ~n9402;
  assign n9404 = ~n9400 & n9403;
  assign n9405 = ~n6397 & n9404;
  assign n9406 = ~n4204 & n9404;
  assign n9407 = ~n9405 & ~n9406;
  assign n9408 =  a[14]  & ~n9407;
  assign n9409 = ~ a[14]  & n9407;
  assign n9410 = ~n9408 & ~n9409;
  assign n9411 = n9399 & ~n9410;
  assign n9412 = n8957 & n9285;
  assign n9413 = ~n9286 & ~n9412;
  assign n9414 = ~n958 & n7101;
  assign n9415 = ~n1178 & n6402;
  assign n9416 = ~n1060 & n6951;
  assign n9417 = ~n9415 & ~n9416;
  assign n9418 = ~n9414 & n9417;
  assign n9419 = ~n6397 & n9418;
  assign n9420 = ~n4633 & n9418;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 =  a[14]  & ~n9421;
  assign n9423 = ~ a[14]  & n9421;
  assign n9424 = ~n9422 & ~n9423;
  assign n9425 = n9413 & ~n9424;
  assign n9426 = n8975 & n9283;
  assign n9427 = ~n9284 & ~n9426;
  assign n9428 = ~n1060 & n7101;
  assign n9429 = ~n1235 & n6402;
  assign n9430 = ~n1178 & n6951;
  assign n9431 = ~n9429 & ~n9430;
  assign n9432 = ~n9428 & n9431;
  assign n9433 = ~n6397 & n9432;
  assign n9434 = ~n4429 & n9432;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 =  a[14]  & ~n9435;
  assign n9437 = ~ a[14]  & n9435;
  assign n9438 = ~n9436 & ~n9437;
  assign n9439 = n9427 & ~n9438;
  assign n9440 = n8993 & n9281;
  assign n9441 = ~n9282 & ~n9440;
  assign n9442 = ~n1178 & n7101;
  assign n9443 = ~n1364 & n6402;
  assign n9444 = ~n1235 & n6951;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = ~n9442 & n9445;
  assign n9447 = ~n6397 & n9446;
  assign n9448 = ~n4861 & n9446;
  assign n9449 = ~n9447 & ~n9448;
  assign n9450 =  a[14]  & ~n9449;
  assign n9451 = ~ a[14]  & n9449;
  assign n9452 = ~n9450 & ~n9451;
  assign n9453 = n9441 & ~n9452;
  assign n9454 = n9011 & n9279;
  assign n9455 = ~n9280 & ~n9454;
  assign n9456 = ~n1235 & n7101;
  assign n9457 = ~n1472 & n6402;
  assign n9458 = ~n1364 & n6951;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = ~n9456 & n9459;
  assign n9461 = ~n6397 & n9460;
  assign n9462 = ~n4848 & n9460;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 =  a[14]  & ~n9463;
  assign n9465 = ~ a[14]  & n9463;
  assign n9466 = ~n9464 & ~n9465;
  assign n9467 = n9455 & ~n9466;
  assign n9468 = ~n1364 & n7101;
  assign n9469 = ~n1572 & n6402;
  assign n9470 = ~n1472 & n6951;
  assign n9471 = ~n9469 & ~n9470;
  assign n9472 = ~n9468 & n9471;
  assign n9473 = n5114 & n6397;
  assign n9474 = n9472 & ~n9473;
  assign n9475 =  a[14]  & ~n9474;
  assign n9476 = ~n9474 & ~n9475;
  assign n9477 =  a[14]  & ~n9475;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = n9275 & ~n9277;
  assign n9480 = ~n9278 & ~n9479;
  assign n9481 = ~n9478 & n9480;
  assign n9482 = ~n9478 & ~n9481;
  assign n9483 = n9480 & ~n9481;
  assign n9484 = ~n9482 & ~n9483;
  assign n9485 = ~n1472 & n7101;
  assign n9486 = ~n1665 & n6402;
  assign n9487 = ~n1572 & n6951;
  assign n9488 = ~n9486 & ~n9487;
  assign n9489 = ~n9485 & n9488;
  assign n9490 = n5139 & n6397;
  assign n9491 = n9489 & ~n9490;
  assign n9492 =  a[14]  & ~n9491;
  assign n9493 = ~n9491 & ~n9492;
  assign n9494 =  a[14]  & ~n9492;
  assign n9495 = ~n9493 & ~n9494;
  assign n9496 = ~n9270 & ~n9274;
  assign n9497 = ~n9273 & ~n9274;
  assign n9498 = ~n9496 & ~n9497;
  assign n9499 = ~n9495 & ~n9498;
  assign n9500 = ~n9495 & ~n9499;
  assign n9501 = ~n9498 & ~n9499;
  assign n9502 = ~n9500 & ~n9501;
  assign n9503 = n9056 & n9268;
  assign n9504 = ~n9269 & ~n9503;
  assign n9505 = ~n1572 & n7101;
  assign n9506 = ~n1779 & n6402;
  assign n9507 = ~n1665 & n6951;
  assign n9508 = ~n9506 & ~n9507;
  assign n9509 = ~n9505 & n9508;
  assign n9510 = ~n6397 & n9509;
  assign n9511 = ~n5561 & n9509;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 =  a[14]  & ~n9512;
  assign n9514 = ~ a[14]  & n9512;
  assign n9515 = ~n9513 & ~n9514;
  assign n9516 = n9504 & ~n9515;
  assign n9517 = n9074 & n9266;
  assign n9518 = ~n9267 & ~n9517;
  assign n9519 = ~n1665 & n7101;
  assign n9520 = ~n1877 & n6402;
  assign n9521 = ~n1779 & n6951;
  assign n9522 = ~n9520 & ~n9521;
  assign n9523 = ~n9519 & n9522;
  assign n9524 = ~n6397 & n9523;
  assign n9525 = ~n5328 & n9523;
  assign n9526 = ~n9524 & ~n9525;
  assign n9527 =  a[14]  & ~n9526;
  assign n9528 = ~ a[14]  & n9526;
  assign n9529 = ~n9527 & ~n9528;
  assign n9530 = n9518 & ~n9529;
  assign n9531 = n9092 & n9264;
  assign n9532 = ~n9265 & ~n9531;
  assign n9533 = ~n1779 & n7101;
  assign n9534 = ~n1913 & n6402;
  assign n9535 = ~n1877 & n6951;
  assign n9536 = ~n9534 & ~n9535;
  assign n9537 = ~n9533 & n9536;
  assign n9538 = ~n6397 & n9537;
  assign n9539 = ~n5851 & n9537;
  assign n9540 = ~n9538 & ~n9539;
  assign n9541 =  a[14]  & ~n9540;
  assign n9542 = ~ a[14]  & n9540;
  assign n9543 = ~n9541 & ~n9542;
  assign n9544 = n9532 & ~n9543;
  assign n9545 = ~n1877 & n7101;
  assign n9546 = ~n1992 & n6402;
  assign n9547 = ~n1913 & n6951;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = ~n9545 & n9548;
  assign n9550 = n6007 & n6397;
  assign n9551 = n9549 & ~n9550;
  assign n9552 =  a[14]  & ~n9551;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 =  a[14]  & ~n9552;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = n9260 & ~n9262;
  assign n9557 = ~n9263 & ~n9556;
  assign n9558 = ~n9555 & n9557;
  assign n9559 = ~n9555 & ~n9558;
  assign n9560 = n9557 & ~n9558;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = ~n1913 & n7101;
  assign n9563 = ~n2057 & n6402;
  assign n9564 = ~n1992 & n6951;
  assign n9565 = ~n9563 & ~n9564;
  assign n9566 = ~n9562 & n9565;
  assign n9567 = n5834 & n6397;
  assign n9568 = n9566 & ~n9567;
  assign n9569 =  a[14]  & ~n9568;
  assign n9570 = ~n9568 & ~n9569;
  assign n9571 =  a[14]  & ~n9569;
  assign n9572 = ~n9570 & ~n9571;
  assign n9573 = ~n9255 & ~n9259;
  assign n9574 = ~n9258 & ~n9259;
  assign n9575 = ~n9573 & ~n9574;
  assign n9576 = ~n9572 & ~n9575;
  assign n9577 = ~n9572 & ~n9576;
  assign n9578 = ~n9575 & ~n9576;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = ~n1992 & n7101;
  assign n9581 = ~n2152 & n6402;
  assign n9582 = ~n2057 & n6951;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = ~n9580 & n9583;
  assign n9585 = n6143 & n6397;
  assign n9586 = n9584 & ~n9585;
  assign n9587 =  a[14]  & ~n9586;
  assign n9588 = ~n9586 & ~n9587;
  assign n9589 =  a[14]  & ~n9587;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = ~n9250 & ~n9254;
  assign n9592 = ~n9253 & ~n9254;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = ~n9590 & ~n9593;
  assign n9595 = ~n9590 & ~n9594;
  assign n9596 = ~n9593 & ~n9594;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = n9151 & n9248;
  assign n9599 = ~n9249 & ~n9598;
  assign n9600 = ~n2057 & n7101;
  assign n9601 = ~n2189 & n6402;
  assign n9602 = ~n2152 & n6951;
  assign n9603 = ~n9601 & ~n9602;
  assign n9604 = ~n9600 & n9603;
  assign n9605 = ~n6397 & n9604;
  assign n9606 = ~n6479 & n9604;
  assign n9607 = ~n9605 & ~n9606;
  assign n9608 =  a[14]  & ~n9607;
  assign n9609 = ~ a[14]  & n9607;
  assign n9610 = ~n9608 & ~n9609;
  assign n9611 = n9599 & ~n9610;
  assign n9612 = n9244 & ~n9246;
  assign n9613 = ~n9247 & ~n9612;
  assign n9614 = ~n2152 & n7101;
  assign n9615 = ~n2291 & n6402;
  assign n9616 = ~n2189 & n6951;
  assign n9617 = ~n9615 & ~n9616;
  assign n9618 = ~n9614 & n9617;
  assign n9619 = ~n6397 & n9618;
  assign n9620 = ~n6492 & n9618;
  assign n9621 = ~n9619 & ~n9620;
  assign n9622 =  a[14]  & ~n9621;
  assign n9623 = ~ a[14]  & n9621;
  assign n9624 = ~n9622 & ~n9623;
  assign n9625 = n9613 & ~n9624;
  assign n9626 = n9183 & n9242;
  assign n9627 = ~n9243 & ~n9626;
  assign n9628 = ~n2189 & n7101;
  assign n9629 = ~n2388 & n6402;
  assign n9630 = ~n2291 & n6951;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = ~n9628 & n9631;
  assign n9633 = ~n6397 & n9632;
  assign n9634 = ~n6122 & n9632;
  assign n9635 = ~n9633 & ~n9634;
  assign n9636 =  a[14]  & ~n9635;
  assign n9637 = ~ a[14]  & n9635;
  assign n9638 = ~n9636 & ~n9637;
  assign n9639 = n9627 & ~n9638;
  assign n9640 = ~n2291 & n7101;
  assign n9641 = ~n2464 & n6402;
  assign n9642 = ~n2388 & n6951;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = ~n9640 & n9643;
  assign n9645 = n6397 & n6541;
  assign n9646 = n9644 & ~n9645;
  assign n9647 =  a[14]  & ~n9646;
  assign n9648 = ~n9646 & ~n9647;
  assign n9649 =  a[14]  & ~n9647;
  assign n9650 = ~n9648 & ~n9649;
  assign n9651 = n9238 & ~n9240;
  assign n9652 = ~n9241 & ~n9651;
  assign n9653 = ~n9650 & n9652;
  assign n9654 = ~n9650 & ~n9653;
  assign n9655 = n9652 & ~n9653;
  assign n9656 = ~n9654 & ~n9655;
  assign n9657 = ~n9225 & ~n9237;
  assign n9658 = ~n9236 & ~n9237;
  assign n9659 = ~n9657 & ~n9658;
  assign n9660 = ~n2388 & n7101;
  assign n9661 = ~n2533 & n6402;
  assign n9662 = ~n2464 & n6951;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = ~n9660 & n9663;
  assign n9665 = ~n6397 & n9664;
  assign n9666 = ~n6591 & n9664;
  assign n9667 = ~n9665 & ~n9666;
  assign n9668 =  a[14]  & ~n9667;
  assign n9669 = ~ a[14]  & n9667;
  assign n9670 = ~n9668 & ~n9669;
  assign n9671 = ~n9659 & ~n9670;
  assign n9672 = ~n2464 & n7101;
  assign n9673 = ~n2571 & n6402;
  assign n9674 = ~n2533 & n6951;
  assign n9675 = ~n9673 & ~n9674;
  assign n9676 = ~n9672 & n9675;
  assign n9677 = n6397 & n6646;
  assign n9678 = n9676 & ~n9677;
  assign n9679 =  a[14]  & ~n9678;
  assign n9680 = ~n9678 & ~n9679;
  assign n9681 =  a[14]  & ~n9679;
  assign n9682 = ~n9680 & ~n9681;
  assign n9683 = ~n9209 & n9220;
  assign n9684 = ~n9221 & ~n9683;
  assign n9685 = ~n9682 & n9684;
  assign n9686 = ~n9682 & ~n9685;
  assign n9687 = n9684 & ~n9685;
  assign n9688 = ~n9686 & ~n9687;
  assign n9689 = n9206 & ~n9208;
  assign n9690 = ~n9209 & ~n9689;
  assign n9691 = ~n2533 & n7101;
  assign n9692 = ~n2674 & n6402;
  assign n9693 = ~n2571 & n6951;
  assign n9694 = ~n9692 & ~n9693;
  assign n9695 = ~n9691 & n9694;
  assign n9696 = ~n6397 & n9695;
  assign n9697 = ~n6695 & n9695;
  assign n9698 = ~n9696 & ~n9697;
  assign n9699 =  a[14]  & ~n9698;
  assign n9700 = ~ a[14]  & n9698;
  assign n9701 = ~n9699 & ~n9700;
  assign n9702 = n9690 & ~n9701;
  assign n9703 = ~n2829 & n6951;
  assign n9704 = ~n2736 & n7101;
  assign n9705 = ~n9703 & ~n9704;
  assign n9706 = n6397 & ~n7469;
  assign n9707 = n9705 & ~n9706;
  assign n9708 =  a[14]  & ~n9707;
  assign n9709 =  a[14]  & ~n9708;
  assign n9710 = ~n9707 & ~n9708;
  assign n9711 = ~n9709 & ~n9710;
  assign n9712 = ~n2829 & ~n6393;
  assign n9713 =  a[14]  & ~n9712;
  assign n9714 = ~n9711 & n9713;
  assign n9715 = ~n2674 & n7101;
  assign n9716 = ~n2829 & n6402;
  assign n9717 = ~n2736 & n6951;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = ~n9715 & n9718;
  assign n9720 = ~n6397 & n9719;
  assign n9721 = ~n6798 & n9719;
  assign n9722 = ~n9720 & ~n9721;
  assign n9723 =  a[14]  & ~n9722;
  assign n9724 = ~ a[14]  & n9722;
  assign n9725 = ~n9723 & ~n9724;
  assign n9726 = n9714 & ~n9725;
  assign n9727 = n9207 & n9726;
  assign n9728 = n9726 & ~n9727;
  assign n9729 = n9207 & ~n9727;
  assign n9730 = ~n9728 & ~n9729;
  assign n9731 = ~n2571 & n7101;
  assign n9732 = ~n2736 & n6402;
  assign n9733 = ~n2674 & n6951;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = ~n9731 & n9734;
  assign n9736 = n6397 & n6806;
  assign n9737 = n9735 & ~n9736;
  assign n9738 =  a[14]  & ~n9737;
  assign n9739 =  a[14]  & ~n9738;
  assign n9740 = ~n9737 & ~n9738;
  assign n9741 = ~n9739 & ~n9740;
  assign n9742 = ~n9730 & ~n9741;
  assign n9743 = ~n9727 & ~n9742;
  assign n9744 = ~n9690 & n9701;
  assign n9745 = ~n9702 & ~n9744;
  assign n9746 = ~n9743 & n9745;
  assign n9747 = ~n9702 & ~n9746;
  assign n9748 = ~n9688 & ~n9747;
  assign n9749 = ~n9685 & ~n9748;
  assign n9750 = n9659 & n9670;
  assign n9751 = ~n9671 & ~n9750;
  assign n9752 = ~n9749 & n9751;
  assign n9753 = ~n9671 & ~n9752;
  assign n9754 = ~n9656 & ~n9753;
  assign n9755 = ~n9653 & ~n9754;
  assign n9756 = n9627 & ~n9639;
  assign n9757 = ~n9638 & ~n9639;
  assign n9758 = ~n9756 & ~n9757;
  assign n9759 = ~n9755 & ~n9758;
  assign n9760 = ~n9639 & ~n9759;
  assign n9761 = n9613 & ~n9625;
  assign n9762 = ~n9624 & ~n9625;
  assign n9763 = ~n9761 & ~n9762;
  assign n9764 = ~n9760 & ~n9763;
  assign n9765 = ~n9625 & ~n9764;
  assign n9766 = ~n9599 & n9610;
  assign n9767 = ~n9611 & ~n9766;
  assign n9768 = ~n9765 & n9767;
  assign n9769 = ~n9611 & ~n9768;
  assign n9770 = ~n9597 & ~n9769;
  assign n9771 = ~n9594 & ~n9770;
  assign n9772 = ~n9579 & ~n9771;
  assign n9773 = ~n9576 & ~n9772;
  assign n9774 = ~n9561 & ~n9773;
  assign n9775 = ~n9558 & ~n9774;
  assign n9776 = n9532 & ~n9544;
  assign n9777 = ~n9543 & ~n9544;
  assign n9778 = ~n9776 & ~n9777;
  assign n9779 = ~n9775 & ~n9778;
  assign n9780 = ~n9544 & ~n9779;
  assign n9781 = n9518 & ~n9530;
  assign n9782 = ~n9529 & ~n9530;
  assign n9783 = ~n9781 & ~n9782;
  assign n9784 = ~n9780 & ~n9783;
  assign n9785 = ~n9530 & ~n9784;
  assign n9786 = ~n9504 & n9515;
  assign n9787 = ~n9516 & ~n9786;
  assign n9788 = ~n9785 & n9787;
  assign n9789 = ~n9516 & ~n9788;
  assign n9790 = ~n9502 & ~n9789;
  assign n9791 = ~n9499 & ~n9790;
  assign n9792 = ~n9484 & ~n9791;
  assign n9793 = ~n9481 & ~n9792;
  assign n9794 = n9455 & ~n9467;
  assign n9795 = ~n9466 & ~n9467;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = ~n9793 & ~n9796;
  assign n9798 = ~n9467 & ~n9797;
  assign n9799 = n9441 & ~n9453;
  assign n9800 = ~n9452 & ~n9453;
  assign n9801 = ~n9799 & ~n9800;
  assign n9802 = ~n9798 & ~n9801;
  assign n9803 = ~n9453 & ~n9802;
  assign n9804 = n9427 & ~n9439;
  assign n9805 = ~n9438 & ~n9439;
  assign n9806 = ~n9804 & ~n9805;
  assign n9807 = ~n9803 & ~n9806;
  assign n9808 = ~n9439 & ~n9807;
  assign n9809 = n9413 & ~n9425;
  assign n9810 = ~n9424 & ~n9425;
  assign n9811 = ~n9809 & ~n9810;
  assign n9812 = ~n9808 & ~n9811;
  assign n9813 = ~n9425 & ~n9812;
  assign n9814 = n9399 & ~n9411;
  assign n9815 = ~n9410 & ~n9411;
  assign n9816 = ~n9814 & ~n9815;
  assign n9817 = ~n9813 & ~n9816;
  assign n9818 = ~n9411 & ~n9817;
  assign n9819 = n9385 & ~n9397;
  assign n9820 = ~n9396 & ~n9397;
  assign n9821 = ~n9819 & ~n9820;
  assign n9822 = ~n9818 & ~n9821;
  assign n9823 = ~n9397 & ~n9822;
  assign n9824 = n9371 & ~n9383;
  assign n9825 = ~n9382 & ~n9383;
  assign n9826 = ~n9824 & ~n9825;
  assign n9827 = ~n9823 & ~n9826;
  assign n9828 = ~n9383 & ~n9827;
  assign n9829 = n9307 & ~n9309;
  assign n9830 = ~n9310 & ~n9829;
  assign n9831 = ~n9828 & n9830;
  assign n9832 = ~n3605 & n7983;
  assign n9833 = ~n3012 & n7291;
  assign n9834 = ~n3539 & n7632;
  assign n9835 = ~n9833 & ~n9834;
  assign n9836 = ~n9832 & n9835;
  assign n9837 = n4084 & n7294;
  assign n9838 = n9836 & ~n9837;
  assign n9839 =  a[11]  & ~n9838;
  assign n9840 = ~n9838 & ~n9839;
  assign n9841 =  a[11]  & ~n9839;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = n9828 & ~n9830;
  assign n9844 = ~n9831 & ~n9843;
  assign n9845 = ~n9842 & n9844;
  assign n9846 = ~n9831 & ~n9845;
  assign n9847 = ~n9369 & ~n9846;
  assign n9848 = n9369 & n9846;
  assign n9849 = ~n9847 & ~n9848;
  assign n9850 = ~n4045 & n9331;
  assign n9851 = ~n3805 & n8418;
  assign n9852 = ~n3964 & n8860;
  assign n9853 = ~n9851 & ~n9852;
  assign n9854 = ~n9850 & n9853;
  assign n9855 = n4477 & n8421;
  assign n9856 = n9854 & ~n9855;
  assign n9857 =  a[8]  & ~n9856;
  assign n9858 =  a[8]  & ~n9857;
  assign n9859 = ~n9856 & ~n9857;
  assign n9860 = ~n9858 & ~n9859;
  assign n9861 = n9849 & ~n9860;
  assign n9862 = ~n9847 & ~n9861;
  assign n9863 = ~ a[3]  &  a[4] ;
  assign n9864 =  a[3]  & ~ a[4] ;
  assign n9865 = ~n9863 & ~n9864;
  assign n9866 = ~n67 & n70;
  assign n9867 = n9865 & n9866;
  assign n9868 = ~n4515 & n9867;
  assign n9869 = ~n4522 & ~n9868;
  assign n9870 = ~n67 & ~n70;
  assign n9871 = ~n9868 & ~n9870;
  assign n9872 = ~n9869 & ~n9871;
  assign n9873 =  a[5]  & ~n9872;
  assign n9874 = ~ a[5]  & n9872;
  assign n9875 = ~n9873 & ~n9874;
  assign n9876 = ~n9862 & ~n9875;
  assign n9877 = n9330 & ~n9343;
  assign n9878 = ~n9342 & ~n9343;
  assign n9879 = ~n9877 & ~n9878;
  assign n9880 = n9862 & n9875;
  assign n9881 = ~n9876 & ~n9880;
  assign n9882 = ~n9879 & n9881;
  assign n9883 = ~n9876 & ~n9882;
  assign n9884 = ~n9358 & ~n9361;
  assign n9885 = ~n9357 & n9884;
  assign n9886 = ~n9362 & ~n9885;
  assign n9887 = ~n9883 & n9886;
  assign n9888 = ~n9879 & ~n9882;
  assign n9889 = n9881 & ~n9882;
  assign n9890 = ~n9888 & ~n9889;
  assign n9891 = ~n3539 & n7983;
  assign n9892 = ~n392 & n7291;
  assign n9893 = ~n3012 & n7632;
  assign n9894 = ~n9892 & ~n9893;
  assign n9895 = ~n9891 & n9894;
  assign n9896 = n3715 & n7294;
  assign n9897 = n9895 & ~n9896;
  assign n9898 =  a[11]  & ~n9897;
  assign n9899 = ~n9897 & ~n9898;
  assign n9900 =  a[11]  & ~n9898;
  assign n9901 = ~n9899 & ~n9900;
  assign n9902 = ~n9823 & ~n9827;
  assign n9903 = ~n9826 & ~n9827;
  assign n9904 = ~n9902 & ~n9903;
  assign n9905 = ~n9901 & ~n9904;
  assign n9906 = ~n9901 & ~n9905;
  assign n9907 = ~n9904 & ~n9905;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = ~n3012 & n7983;
  assign n9910 = ~n587 & n7291;
  assign n9911 = ~n392 & n7632;
  assign n9912 = ~n9910 & ~n9911;
  assign n9913 = ~n9909 & n9912;
  assign n9914 = n3018 & n7294;
  assign n9915 = n9913 & ~n9914;
  assign n9916 =  a[11]  & ~n9915;
  assign n9917 = ~n9915 & ~n9916;
  assign n9918 =  a[11]  & ~n9916;
  assign n9919 = ~n9917 & ~n9918;
  assign n9920 = ~n9818 & ~n9822;
  assign n9921 = ~n9821 & ~n9822;
  assign n9922 = ~n9920 & ~n9921;
  assign n9923 = ~n9919 & ~n9922;
  assign n9924 = ~n9919 & ~n9923;
  assign n9925 = ~n9922 & ~n9923;
  assign n9926 = ~n9924 & ~n9925;
  assign n9927 = ~n392 & n7983;
  assign n9928 = ~n710 & n7291;
  assign n9929 = ~n587 & n7632;
  assign n9930 = ~n9928 & ~n9929;
  assign n9931 = ~n9927 & n9930;
  assign n9932 = n3347 & n7294;
  assign n9933 = n9931 & ~n9932;
  assign n9934 =  a[11]  & ~n9933;
  assign n9935 = ~n9933 & ~n9934;
  assign n9936 =  a[11]  & ~n9934;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = ~n9813 & ~n9817;
  assign n9939 = ~n9816 & ~n9817;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = ~n9937 & ~n9940;
  assign n9942 = ~n9937 & ~n9941;
  assign n9943 = ~n9940 & ~n9941;
  assign n9944 = ~n9942 & ~n9943;
  assign n9945 = ~n587 & n7983;
  assign n9946 = ~n867 & n7291;
  assign n9947 = ~n710 & n7632;
  assign n9948 = ~n9946 & ~n9947;
  assign n9949 = ~n9945 & n9948;
  assign n9950 = n3331 & n7294;
  assign n9951 = n9949 & ~n9950;
  assign n9952 =  a[11]  & ~n9951;
  assign n9953 = ~n9951 & ~n9952;
  assign n9954 =  a[11]  & ~n9952;
  assign n9955 = ~n9953 & ~n9954;
  assign n9956 = ~n9808 & ~n9812;
  assign n9957 = ~n9811 & ~n9812;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = ~n9955 & ~n9958;
  assign n9960 = ~n9955 & ~n9959;
  assign n9961 = ~n9958 & ~n9959;
  assign n9962 = ~n9960 & ~n9961;
  assign n9963 = ~n710 & n7983;
  assign n9964 = ~n958 & n7291;
  assign n9965 = ~n867 & n7632;
  assign n9966 = ~n9964 & ~n9965;
  assign n9967 = ~n9963 & n9966;
  assign n9968 = n4179 & n7294;
  assign n9969 = n9967 & ~n9968;
  assign n9970 =  a[11]  & ~n9969;
  assign n9971 = ~n9969 & ~n9970;
  assign n9972 =  a[11]  & ~n9970;
  assign n9973 = ~n9971 & ~n9972;
  assign n9974 = ~n9803 & ~n9807;
  assign n9975 = ~n9806 & ~n9807;
  assign n9976 = ~n9974 & ~n9975;
  assign n9977 = ~n9973 & ~n9976;
  assign n9978 = ~n9973 & ~n9977;
  assign n9979 = ~n9976 & ~n9977;
  assign n9980 = ~n9978 & ~n9979;
  assign n9981 = ~n867 & n7983;
  assign n9982 = ~n1060 & n7291;
  assign n9983 = ~n958 & n7632;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = ~n9981 & n9984;
  assign n9986 = n4204 & n7294;
  assign n9987 = n9985 & ~n9986;
  assign n9988 =  a[11]  & ~n9987;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 =  a[11]  & ~n9988;
  assign n9991 = ~n9989 & ~n9990;
  assign n9992 = ~n9798 & ~n9802;
  assign n9993 = ~n9801 & ~n9802;
  assign n9994 = ~n9992 & ~n9993;
  assign n9995 = ~n9991 & ~n9994;
  assign n9996 = ~n9991 & ~n9995;
  assign n9997 = ~n9994 & ~n9995;
  assign n9998 = ~n9996 & ~n9997;
  assign n9999 = ~n958 & n7983;
  assign n10000 = ~n1178 & n7291;
  assign n10001 = ~n1060 & n7632;
  assign n10002 = ~n10000 & ~n10001;
  assign n10003 = ~n9999 & n10002;
  assign n10004 = n4633 & n7294;
  assign n10005 = n10003 & ~n10004;
  assign n10006 =  a[11]  & ~n10005;
  assign n10007 = ~n10005 & ~n10006;
  assign n10008 =  a[11]  & ~n10006;
  assign n10009 = ~n10007 & ~n10008;
  assign n10010 = ~n9793 & ~n9797;
  assign n10011 = ~n9796 & ~n9797;
  assign n10012 = ~n10010 & ~n10011;
  assign n10013 = ~n10009 & ~n10012;
  assign n10014 = ~n10009 & ~n10013;
  assign n10015 = ~n10012 & ~n10013;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = n9484 & n9791;
  assign n10018 = ~n9792 & ~n10017;
  assign n10019 = ~n1060 & n7983;
  assign n10020 = ~n1235 & n7291;
  assign n10021 = ~n1178 & n7632;
  assign n10022 = ~n10020 & ~n10021;
  assign n10023 = ~n10019 & n10022;
  assign n10024 = ~n7294 & n10023;
  assign n10025 = ~n4429 & n10023;
  assign n10026 = ~n10024 & ~n10025;
  assign n10027 =  a[11]  & ~n10026;
  assign n10028 = ~ a[11]  & n10026;
  assign n10029 = ~n10027 & ~n10028;
  assign n10030 = n10018 & ~n10029;
  assign n10031 = n9502 & n9789;
  assign n10032 = ~n9790 & ~n10031;
  assign n10033 = ~n1178 & n7983;
  assign n10034 = ~n1364 & n7291;
  assign n10035 = ~n1235 & n7632;
  assign n10036 = ~n10034 & ~n10035;
  assign n10037 = ~n10033 & n10036;
  assign n10038 = ~n7294 & n10037;
  assign n10039 = ~n4861 & n10037;
  assign n10040 = ~n10038 & ~n10039;
  assign n10041 =  a[11]  & ~n10040;
  assign n10042 = ~ a[11]  & n10040;
  assign n10043 = ~n10041 & ~n10042;
  assign n10044 = n10032 & ~n10043;
  assign n10045 = ~n1235 & n7983;
  assign n10046 = ~n1472 & n7291;
  assign n10047 = ~n1364 & n7632;
  assign n10048 = ~n10046 & ~n10047;
  assign n10049 = ~n10045 & n10048;
  assign n10050 = n4848 & n7294;
  assign n10051 = n10049 & ~n10050;
  assign n10052 =  a[11]  & ~n10051;
  assign n10053 = ~n10051 & ~n10052;
  assign n10054 =  a[11]  & ~n10052;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = n9785 & ~n9787;
  assign n10057 = ~n9788 & ~n10056;
  assign n10058 = ~n10055 & n10057;
  assign n10059 = ~n10055 & ~n10058;
  assign n10060 = n10057 & ~n10058;
  assign n10061 = ~n10059 & ~n10060;
  assign n10062 = ~n1364 & n7983;
  assign n10063 = ~n1572 & n7291;
  assign n10064 = ~n1472 & n7632;
  assign n10065 = ~n10063 & ~n10064;
  assign n10066 = ~n10062 & n10065;
  assign n10067 = n5114 & n7294;
  assign n10068 = n10066 & ~n10067;
  assign n10069 =  a[11]  & ~n10068;
  assign n10070 = ~n10068 & ~n10069;
  assign n10071 =  a[11]  & ~n10069;
  assign n10072 = ~n10070 & ~n10071;
  assign n10073 = ~n9780 & ~n9784;
  assign n10074 = ~n9783 & ~n9784;
  assign n10075 = ~n10073 & ~n10074;
  assign n10076 = ~n10072 & ~n10075;
  assign n10077 = ~n10072 & ~n10076;
  assign n10078 = ~n10075 & ~n10076;
  assign n10079 = ~n10077 & ~n10078;
  assign n10080 = ~n1472 & n7983;
  assign n10081 = ~n1665 & n7291;
  assign n10082 = ~n1572 & n7632;
  assign n10083 = ~n10081 & ~n10082;
  assign n10084 = ~n10080 & n10083;
  assign n10085 = n5139 & n7294;
  assign n10086 = n10084 & ~n10085;
  assign n10087 =  a[11]  & ~n10086;
  assign n10088 = ~n10086 & ~n10087;
  assign n10089 =  a[11]  & ~n10087;
  assign n10090 = ~n10088 & ~n10089;
  assign n10091 = ~n9775 & ~n9779;
  assign n10092 = ~n9778 & ~n9779;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = ~n10090 & ~n10093;
  assign n10095 = ~n10090 & ~n10094;
  assign n10096 = ~n10093 & ~n10094;
  assign n10097 = ~n10095 & ~n10096;
  assign n10098 = n9561 & n9773;
  assign n10099 = ~n9774 & ~n10098;
  assign n10100 = ~n1572 & n7983;
  assign n10101 = ~n1779 & n7291;
  assign n10102 = ~n1665 & n7632;
  assign n10103 = ~n10101 & ~n10102;
  assign n10104 = ~n10100 & n10103;
  assign n10105 = ~n7294 & n10104;
  assign n10106 = ~n5561 & n10104;
  assign n10107 = ~n10105 & ~n10106;
  assign n10108 =  a[11]  & ~n10107;
  assign n10109 = ~ a[11]  & n10107;
  assign n10110 = ~n10108 & ~n10109;
  assign n10111 = n10099 & ~n10110;
  assign n10112 = n9579 & n9771;
  assign n10113 = ~n9772 & ~n10112;
  assign n10114 = ~n1665 & n7983;
  assign n10115 = ~n1877 & n7291;
  assign n10116 = ~n1779 & n7632;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = ~n10114 & n10117;
  assign n10119 = ~n7294 & n10118;
  assign n10120 = ~n5328 & n10118;
  assign n10121 = ~n10119 & ~n10120;
  assign n10122 =  a[11]  & ~n10121;
  assign n10123 = ~ a[11]  & n10121;
  assign n10124 = ~n10122 & ~n10123;
  assign n10125 = n10113 & ~n10124;
  assign n10126 = n9597 & n9769;
  assign n10127 = ~n9770 & ~n10126;
  assign n10128 = ~n1779 & n7983;
  assign n10129 = ~n1913 & n7291;
  assign n10130 = ~n1877 & n7632;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = ~n10128 & n10131;
  assign n10133 = ~n7294 & n10132;
  assign n10134 = ~n5851 & n10132;
  assign n10135 = ~n10133 & ~n10134;
  assign n10136 =  a[11]  & ~n10135;
  assign n10137 = ~ a[11]  & n10135;
  assign n10138 = ~n10136 & ~n10137;
  assign n10139 = n10127 & ~n10138;
  assign n10140 = ~n1877 & n7983;
  assign n10141 = ~n1992 & n7291;
  assign n10142 = ~n1913 & n7632;
  assign n10143 = ~n10141 & ~n10142;
  assign n10144 = ~n10140 & n10143;
  assign n10145 = n6007 & n7294;
  assign n10146 = n10144 & ~n10145;
  assign n10147 =  a[11]  & ~n10146;
  assign n10148 = ~n10146 & ~n10147;
  assign n10149 =  a[11]  & ~n10147;
  assign n10150 = ~n10148 & ~n10149;
  assign n10151 = n9765 & ~n9767;
  assign n10152 = ~n9768 & ~n10151;
  assign n10153 = ~n10150 & n10152;
  assign n10154 = ~n10150 & ~n10153;
  assign n10155 = n10152 & ~n10153;
  assign n10156 = ~n10154 & ~n10155;
  assign n10157 = ~n1913 & n7983;
  assign n10158 = ~n2057 & n7291;
  assign n10159 = ~n1992 & n7632;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = ~n10157 & n10160;
  assign n10162 = n5834 & n7294;
  assign n10163 = n10161 & ~n10162;
  assign n10164 =  a[11]  & ~n10163;
  assign n10165 = ~n10163 & ~n10164;
  assign n10166 =  a[11]  & ~n10164;
  assign n10167 = ~n10165 & ~n10166;
  assign n10168 = ~n9760 & ~n9764;
  assign n10169 = ~n9763 & ~n9764;
  assign n10170 = ~n10168 & ~n10169;
  assign n10171 = ~n10167 & ~n10170;
  assign n10172 = ~n10167 & ~n10171;
  assign n10173 = ~n10170 & ~n10171;
  assign n10174 = ~n10172 & ~n10173;
  assign n10175 = ~n1992 & n7983;
  assign n10176 = ~n2152 & n7291;
  assign n10177 = ~n2057 & n7632;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = ~n10175 & n10178;
  assign n10180 = n6143 & n7294;
  assign n10181 = n10179 & ~n10180;
  assign n10182 =  a[11]  & ~n10181;
  assign n10183 = ~n10181 & ~n10182;
  assign n10184 =  a[11]  & ~n10182;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = ~n9755 & ~n9759;
  assign n10187 = ~n9758 & ~n9759;
  assign n10188 = ~n10186 & ~n10187;
  assign n10189 = ~n10185 & ~n10188;
  assign n10190 = ~n10185 & ~n10189;
  assign n10191 = ~n10188 & ~n10189;
  assign n10192 = ~n10190 & ~n10191;
  assign n10193 = n9656 & n9753;
  assign n10194 = ~n9754 & ~n10193;
  assign n10195 = ~n2057 & n7983;
  assign n10196 = ~n2189 & n7291;
  assign n10197 = ~n2152 & n7632;
  assign n10198 = ~n10196 & ~n10197;
  assign n10199 = ~n10195 & n10198;
  assign n10200 = ~n7294 & n10199;
  assign n10201 = ~n6479 & n10199;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 =  a[11]  & ~n10202;
  assign n10204 = ~ a[11]  & n10202;
  assign n10205 = ~n10203 & ~n10204;
  assign n10206 = n10194 & ~n10205;
  assign n10207 = n9749 & ~n9751;
  assign n10208 = ~n9752 & ~n10207;
  assign n10209 = ~n2152 & n7983;
  assign n10210 = ~n2291 & n7291;
  assign n10211 = ~n2189 & n7632;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = ~n10209 & n10212;
  assign n10214 = ~n7294 & n10213;
  assign n10215 = ~n6492 & n10213;
  assign n10216 = ~n10214 & ~n10215;
  assign n10217 =  a[11]  & ~n10216;
  assign n10218 = ~ a[11]  & n10216;
  assign n10219 = ~n10217 & ~n10218;
  assign n10220 = n10208 & ~n10219;
  assign n10221 = n9688 & n9747;
  assign n10222 = ~n9748 & ~n10221;
  assign n10223 = ~n2189 & n7983;
  assign n10224 = ~n2388 & n7291;
  assign n10225 = ~n2291 & n7632;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = ~n10223 & n10226;
  assign n10228 = ~n7294 & n10227;
  assign n10229 = ~n6122 & n10227;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 =  a[11]  & ~n10230;
  assign n10232 = ~ a[11]  & n10230;
  assign n10233 = ~n10231 & ~n10232;
  assign n10234 = n10222 & ~n10233;
  assign n10235 = ~n2291 & n7983;
  assign n10236 = ~n2464 & n7291;
  assign n10237 = ~n2388 & n7632;
  assign n10238 = ~n10236 & ~n10237;
  assign n10239 = ~n10235 & n10238;
  assign n10240 = n6541 & n7294;
  assign n10241 = n10239 & ~n10240;
  assign n10242 =  a[11]  & ~n10241;
  assign n10243 = ~n10241 & ~n10242;
  assign n10244 =  a[11]  & ~n10242;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = n9743 & ~n9745;
  assign n10247 = ~n9746 & ~n10246;
  assign n10248 = ~n10245 & n10247;
  assign n10249 = ~n10245 & ~n10248;
  assign n10250 = n10247 & ~n10248;
  assign n10251 = ~n10249 & ~n10250;
  assign n10252 = ~n9730 & ~n9742;
  assign n10253 = ~n9741 & ~n9742;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = ~n2388 & n7983;
  assign n10256 = ~n2533 & n7291;
  assign n10257 = ~n2464 & n7632;
  assign n10258 = ~n10256 & ~n10257;
  assign n10259 = ~n10255 & n10258;
  assign n10260 = ~n7294 & n10259;
  assign n10261 = ~n6591 & n10259;
  assign n10262 = ~n10260 & ~n10261;
  assign n10263 =  a[11]  & ~n10262;
  assign n10264 = ~ a[11]  & n10262;
  assign n10265 = ~n10263 & ~n10264;
  assign n10266 = ~n10254 & ~n10265;
  assign n10267 = ~n2464 & n7983;
  assign n10268 = ~n2571 & n7291;
  assign n10269 = ~n2533 & n7632;
  assign n10270 = ~n10268 & ~n10269;
  assign n10271 = ~n10267 & n10270;
  assign n10272 = n6646 & n7294;
  assign n10273 = n10271 & ~n10272;
  assign n10274 =  a[11]  & ~n10273;
  assign n10275 = ~n10273 & ~n10274;
  assign n10276 =  a[11]  & ~n10274;
  assign n10277 = ~n10275 & ~n10276;
  assign n10278 = ~n9714 & n9725;
  assign n10279 = ~n9726 & ~n10278;
  assign n10280 = ~n10277 & n10279;
  assign n10281 = ~n10277 & ~n10280;
  assign n10282 = n10279 & ~n10280;
  assign n10283 = ~n10281 & ~n10282;
  assign n10284 = n9711 & ~n9713;
  assign n10285 = ~n9714 & ~n10284;
  assign n10286 = ~n2533 & n7983;
  assign n10287 = ~n2674 & n7291;
  assign n10288 = ~n2571 & n7632;
  assign n10289 = ~n10287 & ~n10288;
  assign n10290 = ~n10286 & n10289;
  assign n10291 = ~n7294 & n10290;
  assign n10292 = ~n6695 & n10290;
  assign n10293 = ~n10291 & ~n10292;
  assign n10294 =  a[11]  & ~n10293;
  assign n10295 = ~ a[11]  & n10293;
  assign n10296 = ~n10294 & ~n10295;
  assign n10297 = n10285 & ~n10296;
  assign n10298 = ~n2829 & n7632;
  assign n10299 = ~n2736 & n7983;
  assign n10300 = ~n10298 & ~n10299;
  assign n10301 = n7294 & ~n7469;
  assign n10302 = n10300 & ~n10301;
  assign n10303 =  a[11]  & ~n10302;
  assign n10304 =  a[11]  & ~n10303;
  assign n10305 = ~n10302 & ~n10303;
  assign n10306 = ~n10304 & ~n10305;
  assign n10307 = ~n2829 & ~n7289;
  assign n10308 =  a[11]  & ~n10307;
  assign n10309 = ~n10306 & n10308;
  assign n10310 = ~n2674 & n7983;
  assign n10311 = ~n2829 & n7291;
  assign n10312 = ~n2736 & n7632;
  assign n10313 = ~n10311 & ~n10312;
  assign n10314 = ~n10310 & n10313;
  assign n10315 = ~n7294 & n10314;
  assign n10316 = ~n6798 & n10314;
  assign n10317 = ~n10315 & ~n10316;
  assign n10318 =  a[11]  & ~n10317;
  assign n10319 = ~ a[11]  & n10317;
  assign n10320 = ~n10318 & ~n10319;
  assign n10321 = n10309 & ~n10320;
  assign n10322 = n9712 & n10321;
  assign n10323 = n10321 & ~n10322;
  assign n10324 = n9712 & ~n10322;
  assign n10325 = ~n10323 & ~n10324;
  assign n10326 = ~n2571 & n7983;
  assign n10327 = ~n2736 & n7291;
  assign n10328 = ~n2674 & n7632;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = ~n10326 & n10329;
  assign n10331 = n6806 & n7294;
  assign n10332 = n10330 & ~n10331;
  assign n10333 =  a[11]  & ~n10332;
  assign n10334 =  a[11]  & ~n10333;
  assign n10335 = ~n10332 & ~n10333;
  assign n10336 = ~n10334 & ~n10335;
  assign n10337 = ~n10325 & ~n10336;
  assign n10338 = ~n10322 & ~n10337;
  assign n10339 = ~n10285 & n10296;
  assign n10340 = ~n10297 & ~n10339;
  assign n10341 = ~n10338 & n10340;
  assign n10342 = ~n10297 & ~n10341;
  assign n10343 = ~n10283 & ~n10342;
  assign n10344 = ~n10280 & ~n10343;
  assign n10345 = n10254 & n10265;
  assign n10346 = ~n10266 & ~n10345;
  assign n10347 = ~n10344 & n10346;
  assign n10348 = ~n10266 & ~n10347;
  assign n10349 = ~n10251 & ~n10348;
  assign n10350 = ~n10248 & ~n10349;
  assign n10351 = n10222 & ~n10234;
  assign n10352 = ~n10233 & ~n10234;
  assign n10353 = ~n10351 & ~n10352;
  assign n10354 = ~n10350 & ~n10353;
  assign n10355 = ~n10234 & ~n10354;
  assign n10356 = n10208 & ~n10220;
  assign n10357 = ~n10219 & ~n10220;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = ~n10355 & ~n10358;
  assign n10360 = ~n10220 & ~n10359;
  assign n10361 = ~n10194 & n10205;
  assign n10362 = ~n10206 & ~n10361;
  assign n10363 = ~n10360 & n10362;
  assign n10364 = ~n10206 & ~n10363;
  assign n10365 = ~n10192 & ~n10364;
  assign n10366 = ~n10189 & ~n10365;
  assign n10367 = ~n10174 & ~n10366;
  assign n10368 = ~n10171 & ~n10367;
  assign n10369 = ~n10156 & ~n10368;
  assign n10370 = ~n10153 & ~n10369;
  assign n10371 = n10127 & ~n10139;
  assign n10372 = ~n10138 & ~n10139;
  assign n10373 = ~n10371 & ~n10372;
  assign n10374 = ~n10370 & ~n10373;
  assign n10375 = ~n10139 & ~n10374;
  assign n10376 = n10113 & ~n10125;
  assign n10377 = ~n10124 & ~n10125;
  assign n10378 = ~n10376 & ~n10377;
  assign n10379 = ~n10375 & ~n10378;
  assign n10380 = ~n10125 & ~n10379;
  assign n10381 = ~n10099 & n10110;
  assign n10382 = ~n10111 & ~n10381;
  assign n10383 = ~n10380 & n10382;
  assign n10384 = ~n10111 & ~n10383;
  assign n10385 = ~n10097 & ~n10384;
  assign n10386 = ~n10094 & ~n10385;
  assign n10387 = ~n10079 & ~n10386;
  assign n10388 = ~n10076 & ~n10387;
  assign n10389 = ~n10061 & ~n10388;
  assign n10390 = ~n10058 & ~n10389;
  assign n10391 = n10032 & ~n10044;
  assign n10392 = ~n10043 & ~n10044;
  assign n10393 = ~n10391 & ~n10392;
  assign n10394 = ~n10390 & ~n10393;
  assign n10395 = ~n10044 & ~n10394;
  assign n10396 = ~n10018 & n10029;
  assign n10397 = ~n10030 & ~n10396;
  assign n10398 = ~n10395 & n10397;
  assign n10399 = ~n10030 & ~n10398;
  assign n10400 = ~n10016 & ~n10399;
  assign n10401 = ~n10013 & ~n10400;
  assign n10402 = ~n9998 & ~n10401;
  assign n10403 = ~n9995 & ~n10402;
  assign n10404 = ~n9980 & ~n10403;
  assign n10405 = ~n9977 & ~n10404;
  assign n10406 = ~n9962 & ~n10405;
  assign n10407 = ~n9959 & ~n10406;
  assign n10408 = ~n9944 & ~n10407;
  assign n10409 = ~n9941 & ~n10408;
  assign n10410 = ~n9926 & ~n10409;
  assign n10411 = ~n9923 & ~n10410;
  assign n10412 = ~n9908 & ~n10411;
  assign n10413 = ~n9905 & ~n10412;
  assign n10414 = n9842 & ~n9844;
  assign n10415 = ~n9845 & ~n10414;
  assign n10416 = ~n10413 & n10415;
  assign n10417 = ~n3964 & n9331;
  assign n10418 = ~n3456 & n8418;
  assign n10419 = ~n3805 & n8860;
  assign n10420 = ~n10418 & ~n10419;
  assign n10421 = ~n10417 & n10420;
  assign n10422 = n4558 & n8421;
  assign n10423 = n10421 & ~n10422;
  assign n10424 =  a[8]  & ~n10423;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 =  a[8]  & ~n10424;
  assign n10427 = ~n10425 & ~n10426;
  assign n10428 = ~n10413 & ~n10416;
  assign n10429 = n10415 & ~n10416;
  assign n10430 = ~n10428 & ~n10429;
  assign n10431 = ~n10427 & ~n10430;
  assign n10432 = ~n10416 & ~n10431;
  assign n10433 = ~n3877 & n9867;
  assign n10434 = n70 & ~n9865;
  assign n10435 = ~n4515 & n10434;
  assign n10436 = ~n10433 & ~n10435;
  assign n10437 = ~n9870 & n10436;
  assign n10438 = ~n4609 & n10436;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 =  a[5]  & ~n10439;
  assign n10441 = ~ a[5]  & n10439;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = ~n10432 & ~n10442;
  assign n10444 = n9849 & ~n9861;
  assign n10445 = ~n9860 & ~n9861;
  assign n10446 = ~n10444 & ~n10445;
  assign n10447 = n10432 & n10442;
  assign n10448 = ~n10443 & ~n10447;
  assign n10449 = ~n10446 & n10448;
  assign n10450 = ~n10443 & ~n10449;
  assign n10451 = ~n9890 & ~n10450;
  assign n10452 = n9890 & n10450;
  assign n10453 = ~n10451 & ~n10452;
  assign n10454 = n9908 & n10411;
  assign n10455 = ~n10412 & ~n10454;
  assign n10456 = ~n3805 & n9331;
  assign n10457 = ~n3605 & n8418;
  assign n10458 = ~n3456 & n8860;
  assign n10459 = ~n10457 & ~n10458;
  assign n10460 = ~n10456 & n10459;
  assign n10461 = ~n8421 & n10460;
  assign n10462 = ~n3818 & n10460;
  assign n10463 = ~n10461 & ~n10462;
  assign n10464 =  a[8]  & ~n10463;
  assign n10465 = ~ a[8]  & n10463;
  assign n10466 = ~n10464 & ~n10465;
  assign n10467 = n10455 & ~n10466;
  assign n10468 = n9926 & n10409;
  assign n10469 = ~n10410 & ~n10468;
  assign n10470 = ~n3456 & n9331;
  assign n10471 = ~n3539 & n8418;
  assign n10472 = ~n3605 & n8860;
  assign n10473 = ~n10471 & ~n10472;
  assign n10474 = ~n10470 & n10473;
  assign n10475 = ~n8421 & n10474;
  assign n10476 = ~n3627 & n10474;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 =  a[8]  & ~n10477;
  assign n10479 = ~ a[8]  & n10477;
  assign n10480 = ~n10478 & ~n10479;
  assign n10481 = n10469 & ~n10480;
  assign n10482 = n9944 & n10407;
  assign n10483 = ~n10408 & ~n10482;
  assign n10484 = ~n3605 & n9331;
  assign n10485 = ~n3012 & n8418;
  assign n10486 = ~n3539 & n8860;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = ~n10484 & n10487;
  assign n10489 = ~n8421 & n10488;
  assign n10490 = ~n4084 & n10488;
  assign n10491 = ~n10489 & ~n10490;
  assign n10492 =  a[8]  & ~n10491;
  assign n10493 = ~ a[8]  & n10491;
  assign n10494 = ~n10492 & ~n10493;
  assign n10495 = n10483 & ~n10494;
  assign n10496 = n9962 & n10405;
  assign n10497 = ~n10406 & ~n10496;
  assign n10498 = ~n3539 & n9331;
  assign n10499 = ~n392 & n8418;
  assign n10500 = ~n3012 & n8860;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = ~n10498 & n10501;
  assign n10503 = ~n8421 & n10502;
  assign n10504 = ~n3715 & n10502;
  assign n10505 = ~n10503 & ~n10504;
  assign n10506 =  a[8]  & ~n10505;
  assign n10507 = ~ a[8]  & n10505;
  assign n10508 = ~n10506 & ~n10507;
  assign n10509 = n10497 & ~n10508;
  assign n10510 = n9980 & n10403;
  assign n10511 = ~n10404 & ~n10510;
  assign n10512 = ~n3012 & n9331;
  assign n10513 = ~n587 & n8418;
  assign n10514 = ~n392 & n8860;
  assign n10515 = ~n10513 & ~n10514;
  assign n10516 = ~n10512 & n10515;
  assign n10517 = ~n8421 & n10516;
  assign n10518 = ~n3018 & n10516;
  assign n10519 = ~n10517 & ~n10518;
  assign n10520 =  a[8]  & ~n10519;
  assign n10521 = ~ a[8]  & n10519;
  assign n10522 = ~n10520 & ~n10521;
  assign n10523 = n10511 & ~n10522;
  assign n10524 = n9998 & n10401;
  assign n10525 = ~n10402 & ~n10524;
  assign n10526 = ~n392 & n9331;
  assign n10527 = ~n710 & n8418;
  assign n10528 = ~n587 & n8860;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = ~n10526 & n10529;
  assign n10531 = ~n8421 & n10530;
  assign n10532 = ~n3347 & n10530;
  assign n10533 = ~n10531 & ~n10532;
  assign n10534 =  a[8]  & ~n10533;
  assign n10535 = ~ a[8]  & n10533;
  assign n10536 = ~n10534 & ~n10535;
  assign n10537 = n10525 & ~n10536;
  assign n10538 = n10016 & n10399;
  assign n10539 = ~n10400 & ~n10538;
  assign n10540 = ~n587 & n9331;
  assign n10541 = ~n867 & n8418;
  assign n10542 = ~n710 & n8860;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = ~n10540 & n10543;
  assign n10545 = ~n8421 & n10544;
  assign n10546 = ~n3331 & n10544;
  assign n10547 = ~n10545 & ~n10546;
  assign n10548 =  a[8]  & ~n10547;
  assign n10549 = ~ a[8]  & n10547;
  assign n10550 = ~n10548 & ~n10549;
  assign n10551 = n10539 & ~n10550;
  assign n10552 = ~n710 & n9331;
  assign n10553 = ~n958 & n8418;
  assign n10554 = ~n867 & n8860;
  assign n10555 = ~n10553 & ~n10554;
  assign n10556 = ~n10552 & n10555;
  assign n10557 = n4179 & n8421;
  assign n10558 = n10556 & ~n10557;
  assign n10559 =  a[8]  & ~n10558;
  assign n10560 = ~n10558 & ~n10559;
  assign n10561 =  a[8]  & ~n10559;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = n10395 & ~n10397;
  assign n10564 = ~n10398 & ~n10563;
  assign n10565 = ~n10562 & n10564;
  assign n10566 = ~n10562 & ~n10565;
  assign n10567 = n10564 & ~n10565;
  assign n10568 = ~n10566 & ~n10567;
  assign n10569 = ~n867 & n9331;
  assign n10570 = ~n1060 & n8418;
  assign n10571 = ~n958 & n8860;
  assign n10572 = ~n10570 & ~n10571;
  assign n10573 = ~n10569 & n10572;
  assign n10574 = n4204 & n8421;
  assign n10575 = n10573 & ~n10574;
  assign n10576 =  a[8]  & ~n10575;
  assign n10577 = ~n10575 & ~n10576;
  assign n10578 =  a[8]  & ~n10576;
  assign n10579 = ~n10577 & ~n10578;
  assign n10580 = ~n10390 & ~n10394;
  assign n10581 = ~n10393 & ~n10394;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = ~n10579 & ~n10582;
  assign n10584 = ~n10579 & ~n10583;
  assign n10585 = ~n10582 & ~n10583;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = n10061 & n10388;
  assign n10588 = ~n10389 & ~n10587;
  assign n10589 = ~n958 & n9331;
  assign n10590 = ~n1178 & n8418;
  assign n10591 = ~n1060 & n8860;
  assign n10592 = ~n10590 & ~n10591;
  assign n10593 = ~n10589 & n10592;
  assign n10594 = ~n8421 & n10593;
  assign n10595 = ~n4633 & n10593;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 =  a[8]  & ~n10596;
  assign n10598 = ~ a[8]  & n10596;
  assign n10599 = ~n10597 & ~n10598;
  assign n10600 = n10588 & ~n10599;
  assign n10601 = n10079 & n10386;
  assign n10602 = ~n10387 & ~n10601;
  assign n10603 = ~n1060 & n9331;
  assign n10604 = ~n1235 & n8418;
  assign n10605 = ~n1178 & n8860;
  assign n10606 = ~n10604 & ~n10605;
  assign n10607 = ~n10603 & n10606;
  assign n10608 = ~n8421 & n10607;
  assign n10609 = ~n4429 & n10607;
  assign n10610 = ~n10608 & ~n10609;
  assign n10611 =  a[8]  & ~n10610;
  assign n10612 = ~ a[8]  & n10610;
  assign n10613 = ~n10611 & ~n10612;
  assign n10614 = n10602 & ~n10613;
  assign n10615 = n10097 & n10384;
  assign n10616 = ~n10385 & ~n10615;
  assign n10617 = ~n1178 & n9331;
  assign n10618 = ~n1364 & n8418;
  assign n10619 = ~n1235 & n8860;
  assign n10620 = ~n10618 & ~n10619;
  assign n10621 = ~n10617 & n10620;
  assign n10622 = ~n8421 & n10621;
  assign n10623 = ~n4861 & n10621;
  assign n10624 = ~n10622 & ~n10623;
  assign n10625 =  a[8]  & ~n10624;
  assign n10626 = ~ a[8]  & n10624;
  assign n10627 = ~n10625 & ~n10626;
  assign n10628 = n10616 & ~n10627;
  assign n10629 = ~n1235 & n9331;
  assign n10630 = ~n1472 & n8418;
  assign n10631 = ~n1364 & n8860;
  assign n10632 = ~n10630 & ~n10631;
  assign n10633 = ~n10629 & n10632;
  assign n10634 = n4848 & n8421;
  assign n10635 = n10633 & ~n10634;
  assign n10636 =  a[8]  & ~n10635;
  assign n10637 = ~n10635 & ~n10636;
  assign n10638 =  a[8]  & ~n10636;
  assign n10639 = ~n10637 & ~n10638;
  assign n10640 = n10380 & ~n10382;
  assign n10641 = ~n10383 & ~n10640;
  assign n10642 = ~n10639 & n10641;
  assign n10643 = ~n10639 & ~n10642;
  assign n10644 = n10641 & ~n10642;
  assign n10645 = ~n10643 & ~n10644;
  assign n10646 = ~n1364 & n9331;
  assign n10647 = ~n1572 & n8418;
  assign n10648 = ~n1472 & n8860;
  assign n10649 = ~n10647 & ~n10648;
  assign n10650 = ~n10646 & n10649;
  assign n10651 = n5114 & n8421;
  assign n10652 = n10650 & ~n10651;
  assign n10653 =  a[8]  & ~n10652;
  assign n10654 = ~n10652 & ~n10653;
  assign n10655 =  a[8]  & ~n10653;
  assign n10656 = ~n10654 & ~n10655;
  assign n10657 = ~n10375 & ~n10379;
  assign n10658 = ~n10378 & ~n10379;
  assign n10659 = ~n10657 & ~n10658;
  assign n10660 = ~n10656 & ~n10659;
  assign n10661 = ~n10656 & ~n10660;
  assign n10662 = ~n10659 & ~n10660;
  assign n10663 = ~n10661 & ~n10662;
  assign n10664 = ~n1472 & n9331;
  assign n10665 = ~n1665 & n8418;
  assign n10666 = ~n1572 & n8860;
  assign n10667 = ~n10665 & ~n10666;
  assign n10668 = ~n10664 & n10667;
  assign n10669 = n5139 & n8421;
  assign n10670 = n10668 & ~n10669;
  assign n10671 =  a[8]  & ~n10670;
  assign n10672 = ~n10670 & ~n10671;
  assign n10673 =  a[8]  & ~n10671;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = ~n10370 & ~n10374;
  assign n10676 = ~n10373 & ~n10374;
  assign n10677 = ~n10675 & ~n10676;
  assign n10678 = ~n10674 & ~n10677;
  assign n10679 = ~n10674 & ~n10678;
  assign n10680 = ~n10677 & ~n10678;
  assign n10681 = ~n10679 & ~n10680;
  assign n10682 = n10156 & n10368;
  assign n10683 = ~n10369 & ~n10682;
  assign n10684 = ~n1572 & n9331;
  assign n10685 = ~n1779 & n8418;
  assign n10686 = ~n1665 & n8860;
  assign n10687 = ~n10685 & ~n10686;
  assign n10688 = ~n10684 & n10687;
  assign n10689 = ~n8421 & n10688;
  assign n10690 = ~n5561 & n10688;
  assign n10691 = ~n10689 & ~n10690;
  assign n10692 =  a[8]  & ~n10691;
  assign n10693 = ~ a[8]  & n10691;
  assign n10694 = ~n10692 & ~n10693;
  assign n10695 = n10683 & ~n10694;
  assign n10696 = n10174 & n10366;
  assign n10697 = ~n10367 & ~n10696;
  assign n10698 = ~n1665 & n9331;
  assign n10699 = ~n1877 & n8418;
  assign n10700 = ~n1779 & n8860;
  assign n10701 = ~n10699 & ~n10700;
  assign n10702 = ~n10698 & n10701;
  assign n10703 = ~n8421 & n10702;
  assign n10704 = ~n5328 & n10702;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 =  a[8]  & ~n10705;
  assign n10707 = ~ a[8]  & n10705;
  assign n10708 = ~n10706 & ~n10707;
  assign n10709 = n10697 & ~n10708;
  assign n10710 = n10192 & n10364;
  assign n10711 = ~n10365 & ~n10710;
  assign n10712 = ~n1779 & n9331;
  assign n10713 = ~n1913 & n8418;
  assign n10714 = ~n1877 & n8860;
  assign n10715 = ~n10713 & ~n10714;
  assign n10716 = ~n10712 & n10715;
  assign n10717 = ~n8421 & n10716;
  assign n10718 = ~n5851 & n10716;
  assign n10719 = ~n10717 & ~n10718;
  assign n10720 =  a[8]  & ~n10719;
  assign n10721 = ~ a[8]  & n10719;
  assign n10722 = ~n10720 & ~n10721;
  assign n10723 = n10711 & ~n10722;
  assign n10724 = ~n1877 & n9331;
  assign n10725 = ~n1992 & n8418;
  assign n10726 = ~n1913 & n8860;
  assign n10727 = ~n10725 & ~n10726;
  assign n10728 = ~n10724 & n10727;
  assign n10729 = n6007 & n8421;
  assign n10730 = n10728 & ~n10729;
  assign n10731 =  a[8]  & ~n10730;
  assign n10732 = ~n10730 & ~n10731;
  assign n10733 =  a[8]  & ~n10731;
  assign n10734 = ~n10732 & ~n10733;
  assign n10735 = n10360 & ~n10362;
  assign n10736 = ~n10363 & ~n10735;
  assign n10737 = ~n10734 & n10736;
  assign n10738 = ~n10734 & ~n10737;
  assign n10739 = n10736 & ~n10737;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = ~n1913 & n9331;
  assign n10742 = ~n2057 & n8418;
  assign n10743 = ~n1992 & n8860;
  assign n10744 = ~n10742 & ~n10743;
  assign n10745 = ~n10741 & n10744;
  assign n10746 = n5834 & n8421;
  assign n10747 = n10745 & ~n10746;
  assign n10748 =  a[8]  & ~n10747;
  assign n10749 = ~n10747 & ~n10748;
  assign n10750 =  a[8]  & ~n10748;
  assign n10751 = ~n10749 & ~n10750;
  assign n10752 = ~n10355 & ~n10359;
  assign n10753 = ~n10358 & ~n10359;
  assign n10754 = ~n10752 & ~n10753;
  assign n10755 = ~n10751 & ~n10754;
  assign n10756 = ~n10751 & ~n10755;
  assign n10757 = ~n10754 & ~n10755;
  assign n10758 = ~n10756 & ~n10757;
  assign n10759 = ~n1992 & n9331;
  assign n10760 = ~n2152 & n8418;
  assign n10761 = ~n2057 & n8860;
  assign n10762 = ~n10760 & ~n10761;
  assign n10763 = ~n10759 & n10762;
  assign n10764 = n6143 & n8421;
  assign n10765 = n10763 & ~n10764;
  assign n10766 =  a[8]  & ~n10765;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 =  a[8]  & ~n10766;
  assign n10769 = ~n10767 & ~n10768;
  assign n10770 = ~n10350 & ~n10354;
  assign n10771 = ~n10353 & ~n10354;
  assign n10772 = ~n10770 & ~n10771;
  assign n10773 = ~n10769 & ~n10772;
  assign n10774 = ~n10769 & ~n10773;
  assign n10775 = ~n10772 & ~n10773;
  assign n10776 = ~n10774 & ~n10775;
  assign n10777 = n10251 & n10348;
  assign n10778 = ~n10349 & ~n10777;
  assign n10779 = ~n2057 & n9331;
  assign n10780 = ~n2189 & n8418;
  assign n10781 = ~n2152 & n8860;
  assign n10782 = ~n10780 & ~n10781;
  assign n10783 = ~n10779 & n10782;
  assign n10784 = ~n8421 & n10783;
  assign n10785 = ~n6479 & n10783;
  assign n10786 = ~n10784 & ~n10785;
  assign n10787 =  a[8]  & ~n10786;
  assign n10788 = ~ a[8]  & n10786;
  assign n10789 = ~n10787 & ~n10788;
  assign n10790 = n10778 & ~n10789;
  assign n10791 = n10344 & ~n10346;
  assign n10792 = ~n10347 & ~n10791;
  assign n10793 = ~n2152 & n9331;
  assign n10794 = ~n2291 & n8418;
  assign n10795 = ~n2189 & n8860;
  assign n10796 = ~n10794 & ~n10795;
  assign n10797 = ~n10793 & n10796;
  assign n10798 = ~n8421 & n10797;
  assign n10799 = ~n6492 & n10797;
  assign n10800 = ~n10798 & ~n10799;
  assign n10801 =  a[8]  & ~n10800;
  assign n10802 = ~ a[8]  & n10800;
  assign n10803 = ~n10801 & ~n10802;
  assign n10804 = n10792 & ~n10803;
  assign n10805 = n10283 & n10342;
  assign n10806 = ~n10343 & ~n10805;
  assign n10807 = ~n2189 & n9331;
  assign n10808 = ~n2388 & n8418;
  assign n10809 = ~n2291 & n8860;
  assign n10810 = ~n10808 & ~n10809;
  assign n10811 = ~n10807 & n10810;
  assign n10812 = ~n8421 & n10811;
  assign n10813 = ~n6122 & n10811;
  assign n10814 = ~n10812 & ~n10813;
  assign n10815 =  a[8]  & ~n10814;
  assign n10816 = ~ a[8]  & n10814;
  assign n10817 = ~n10815 & ~n10816;
  assign n10818 = n10806 & ~n10817;
  assign n10819 = ~n2291 & n9331;
  assign n10820 = ~n2464 & n8418;
  assign n10821 = ~n2388 & n8860;
  assign n10822 = ~n10820 & ~n10821;
  assign n10823 = ~n10819 & n10822;
  assign n10824 = n6541 & n8421;
  assign n10825 = n10823 & ~n10824;
  assign n10826 =  a[8]  & ~n10825;
  assign n10827 = ~n10825 & ~n10826;
  assign n10828 =  a[8]  & ~n10826;
  assign n10829 = ~n10827 & ~n10828;
  assign n10830 = n10338 & ~n10340;
  assign n10831 = ~n10341 & ~n10830;
  assign n10832 = ~n10829 & n10831;
  assign n10833 = ~n10829 & ~n10832;
  assign n10834 = n10831 & ~n10832;
  assign n10835 = ~n10833 & ~n10834;
  assign n10836 = ~n10325 & ~n10337;
  assign n10837 = ~n10336 & ~n10337;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = ~n2388 & n9331;
  assign n10840 = ~n2533 & n8418;
  assign n10841 = ~n2464 & n8860;
  assign n10842 = ~n10840 & ~n10841;
  assign n10843 = ~n10839 & n10842;
  assign n10844 = ~n8421 & n10843;
  assign n10845 = ~n6591 & n10843;
  assign n10846 = ~n10844 & ~n10845;
  assign n10847 =  a[8]  & ~n10846;
  assign n10848 = ~ a[8]  & n10846;
  assign n10849 = ~n10847 & ~n10848;
  assign n10850 = ~n10838 & ~n10849;
  assign n10851 = ~n2464 & n9331;
  assign n10852 = ~n2571 & n8418;
  assign n10853 = ~n2533 & n8860;
  assign n10854 = ~n10852 & ~n10853;
  assign n10855 = ~n10851 & n10854;
  assign n10856 = n6646 & n8421;
  assign n10857 = n10855 & ~n10856;
  assign n10858 =  a[8]  & ~n10857;
  assign n10859 = ~n10857 & ~n10858;
  assign n10860 =  a[8]  & ~n10858;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = ~n10309 & n10320;
  assign n10863 = ~n10321 & ~n10862;
  assign n10864 = ~n10861 & n10863;
  assign n10865 = ~n10861 & ~n10864;
  assign n10866 = n10863 & ~n10864;
  assign n10867 = ~n10865 & ~n10866;
  assign n10868 = n10306 & ~n10308;
  assign n10869 = ~n10309 & ~n10868;
  assign n10870 = ~n2533 & n9331;
  assign n10871 = ~n2674 & n8418;
  assign n10872 = ~n2571 & n8860;
  assign n10873 = ~n10871 & ~n10872;
  assign n10874 = ~n10870 & n10873;
  assign n10875 = ~n8421 & n10874;
  assign n10876 = ~n6695 & n10874;
  assign n10877 = ~n10875 & ~n10876;
  assign n10878 =  a[8]  & ~n10877;
  assign n10879 = ~ a[8]  & n10877;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = n10869 & ~n10880;
  assign n10882 = ~n2829 & n8860;
  assign n10883 = ~n2736 & n9331;
  assign n10884 = ~n10882 & ~n10883;
  assign n10885 = ~n7469 & n8421;
  assign n10886 = n10884 & ~n10885;
  assign n10887 =  a[8]  & ~n10886;
  assign n10888 =  a[8]  & ~n10887;
  assign n10889 = ~n10886 & ~n10887;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = ~n2829 & ~n8416;
  assign n10892 =  a[8]  & ~n10891;
  assign n10893 = ~n10890 & n10892;
  assign n10894 = ~n2674 & n9331;
  assign n10895 = ~n2829 & n8418;
  assign n10896 = ~n2736 & n8860;
  assign n10897 = ~n10895 & ~n10896;
  assign n10898 = ~n10894 & n10897;
  assign n10899 = ~n8421 & n10898;
  assign n10900 = ~n6798 & n10898;
  assign n10901 = ~n10899 & ~n10900;
  assign n10902 =  a[8]  & ~n10901;
  assign n10903 = ~ a[8]  & n10901;
  assign n10904 = ~n10902 & ~n10903;
  assign n10905 = n10893 & ~n10904;
  assign n10906 = n10307 & n10905;
  assign n10907 = n10905 & ~n10906;
  assign n10908 = n10307 & ~n10906;
  assign n10909 = ~n10907 & ~n10908;
  assign n10910 = ~n2571 & n9331;
  assign n10911 = ~n2736 & n8418;
  assign n10912 = ~n2674 & n8860;
  assign n10913 = ~n10911 & ~n10912;
  assign n10914 = ~n10910 & n10913;
  assign n10915 = n6806 & n8421;
  assign n10916 = n10914 & ~n10915;
  assign n10917 =  a[8]  & ~n10916;
  assign n10918 =  a[8]  & ~n10917;
  assign n10919 = ~n10916 & ~n10917;
  assign n10920 = ~n10918 & ~n10919;
  assign n10921 = ~n10909 & ~n10920;
  assign n10922 = ~n10906 & ~n10921;
  assign n10923 = ~n10869 & n10880;
  assign n10924 = ~n10881 & ~n10923;
  assign n10925 = ~n10922 & n10924;
  assign n10926 = ~n10881 & ~n10925;
  assign n10927 = ~n10867 & ~n10926;
  assign n10928 = ~n10864 & ~n10927;
  assign n10929 = n10838 & n10849;
  assign n10930 = ~n10850 & ~n10929;
  assign n10931 = ~n10928 & n10930;
  assign n10932 = ~n10850 & ~n10931;
  assign n10933 = ~n10835 & ~n10932;
  assign n10934 = ~n10832 & ~n10933;
  assign n10935 = n10806 & ~n10818;
  assign n10936 = ~n10817 & ~n10818;
  assign n10937 = ~n10935 & ~n10936;
  assign n10938 = ~n10934 & ~n10937;
  assign n10939 = ~n10818 & ~n10938;
  assign n10940 = n10792 & ~n10804;
  assign n10941 = ~n10803 & ~n10804;
  assign n10942 = ~n10940 & ~n10941;
  assign n10943 = ~n10939 & ~n10942;
  assign n10944 = ~n10804 & ~n10943;
  assign n10945 = ~n10778 & n10789;
  assign n10946 = ~n10790 & ~n10945;
  assign n10947 = ~n10944 & n10946;
  assign n10948 = ~n10790 & ~n10947;
  assign n10949 = ~n10776 & ~n10948;
  assign n10950 = ~n10773 & ~n10949;
  assign n10951 = ~n10758 & ~n10950;
  assign n10952 = ~n10755 & ~n10951;
  assign n10953 = ~n10740 & ~n10952;
  assign n10954 = ~n10737 & ~n10953;
  assign n10955 = n10711 & ~n10723;
  assign n10956 = ~n10722 & ~n10723;
  assign n10957 = ~n10955 & ~n10956;
  assign n10958 = ~n10954 & ~n10957;
  assign n10959 = ~n10723 & ~n10958;
  assign n10960 = n10697 & ~n10709;
  assign n10961 = ~n10708 & ~n10709;
  assign n10962 = ~n10960 & ~n10961;
  assign n10963 = ~n10959 & ~n10962;
  assign n10964 = ~n10709 & ~n10963;
  assign n10965 = ~n10683 & n10694;
  assign n10966 = ~n10695 & ~n10965;
  assign n10967 = ~n10964 & n10966;
  assign n10968 = ~n10695 & ~n10967;
  assign n10969 = ~n10681 & ~n10968;
  assign n10970 = ~n10678 & ~n10969;
  assign n10971 = ~n10663 & ~n10970;
  assign n10972 = ~n10660 & ~n10971;
  assign n10973 = ~n10645 & ~n10972;
  assign n10974 = ~n10642 & ~n10973;
  assign n10975 = n10616 & ~n10628;
  assign n10976 = ~n10627 & ~n10628;
  assign n10977 = ~n10975 & ~n10976;
  assign n10978 = ~n10974 & ~n10977;
  assign n10979 = ~n10628 & ~n10978;
  assign n10980 = n10602 & ~n10614;
  assign n10981 = ~n10613 & ~n10614;
  assign n10982 = ~n10980 & ~n10981;
  assign n10983 = ~n10979 & ~n10982;
  assign n10984 = ~n10614 & ~n10983;
  assign n10985 = ~n10588 & n10599;
  assign n10986 = ~n10600 & ~n10985;
  assign n10987 = ~n10984 & n10986;
  assign n10988 = ~n10600 & ~n10987;
  assign n10989 = ~n10586 & ~n10988;
  assign n10990 = ~n10583 & ~n10989;
  assign n10991 = ~n10568 & ~n10990;
  assign n10992 = ~n10565 & ~n10991;
  assign n10993 = n10539 & ~n10551;
  assign n10994 = ~n10550 & ~n10551;
  assign n10995 = ~n10993 & ~n10994;
  assign n10996 = ~n10992 & ~n10995;
  assign n10997 = ~n10551 & ~n10996;
  assign n10998 = n10525 & ~n10537;
  assign n10999 = ~n10536 & ~n10537;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = ~n10997 & ~n11000;
  assign n11002 = ~n10537 & ~n11001;
  assign n11003 = n10511 & ~n10523;
  assign n11004 = ~n10522 & ~n10523;
  assign n11005 = ~n11003 & ~n11004;
  assign n11006 = ~n11002 & ~n11005;
  assign n11007 = ~n10523 & ~n11006;
  assign n11008 = n10497 & ~n10509;
  assign n11009 = ~n10508 & ~n10509;
  assign n11010 = ~n11008 & ~n11009;
  assign n11011 = ~n11007 & ~n11010;
  assign n11012 = ~n10509 & ~n11011;
  assign n11013 = n10483 & ~n10495;
  assign n11014 = ~n10494 & ~n10495;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = ~n11012 & ~n11015;
  assign n11017 = ~n10495 & ~n11016;
  assign n11018 = n10469 & ~n10481;
  assign n11019 = ~n10480 & ~n10481;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = ~n11017 & ~n11020;
  assign n11022 = ~n10481 & ~n11021;
  assign n11023 = n10455 & ~n10467;
  assign n11024 = ~n10466 & ~n10467;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = ~n11022 & ~n11025;
  assign n11027 = ~n10467 & ~n11026;
  assign n11028 = n10427 & ~n10429;
  assign n11029 = ~n10428 & n11028;
  assign n11030 = ~n10431 & ~n11029;
  assign n11031 = ~n11027 & n11030;
  assign n11032 = n71 & ~n4515;
  assign n11033 = ~n4045 & n9867;
  assign n11034 = ~n3877 & n10434;
  assign n11035 = ~n11033 & ~n11034;
  assign n11036 = ~n11032 & n11035;
  assign n11037 = n4715 & n9870;
  assign n11038 = n11036 & ~n11037;
  assign n11039 =  a[5]  & ~n11038;
  assign n11040 = ~n11038 & ~n11039;
  assign n11041 =  a[5]  & ~n11039;
  assign n11042 = ~n11040 & ~n11041;
  assign n11043 = ~n11027 & ~n11031;
  assign n11044 = n11030 & ~n11031;
  assign n11045 = ~n11043 & ~n11044;
  assign n11046 = ~n11042 & ~n11045;
  assign n11047 = ~n11031 & ~n11046;
  assign n11048 = n10446 & ~n10448;
  assign n11049 = ~n10449 & ~n11048;
  assign n11050 = ~n11047 & n11049;
  assign n11051 =  a[1]  & ~ a[2] ;
  assign n11052 = ~ a[1]  &  a[2] ;
  assign n11053 = ~n11051 & ~n11052;
  assign n11054 = ~ a[0]  & ~ a[1] ;
  assign n11055 = ~n11053 & n11054;
  assign n11056 = ~n4515 & n11055;
  assign n11057 =  a[0]  & ~n11053;
  assign n11058 = n4522 & n11057;
  assign n11059 = ~n11056 & ~n11058;
  assign n11060 =  a[2]  & ~n11059;
  assign n11061 = ~n11059 & ~n11060;
  assign n11062 =  a[2]  & ~n11060;
  assign n11063 = ~n11061 & ~n11062;
  assign n11064 = n71 & ~n3877;
  assign n11065 = ~n3964 & n9867;
  assign n11066 = ~n4045 & n10434;
  assign n11067 = ~n11065 & ~n11066;
  assign n11068 = ~n11064 & n11067;
  assign n11069 = n4067 & n9870;
  assign n11070 = n11068 & ~n11069;
  assign n11071 =  a[5]  & ~n11070;
  assign n11072 =  a[5]  & ~n11071;
  assign n11073 = ~n11070 & ~n11071;
  assign n11074 = ~n11072 & ~n11073;
  assign n11075 = ~n11063 & ~n11074;
  assign n11076 = ~n11063 & ~n11075;
  assign n11077 = ~n11074 & ~n11075;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = ~n11022 & ~n11026;
  assign n11080 = ~n11025 & ~n11026;
  assign n11081 = ~n11079 & ~n11080;
  assign n11082 = ~n11078 & ~n11081;
  assign n11083 = ~n11075 & ~n11082;
  assign n11084 = n11042 & ~n11044;
  assign n11085 = ~n11043 & n11084;
  assign n11086 = ~n11046 & ~n11085;
  assign n11087 = ~n11083 & n11086;
  assign n11088 = ~n11078 & ~n11082;
  assign n11089 = ~n11081 & ~n11082;
  assign n11090 = ~n11088 & ~n11089;
  assign n11091 = n71 & ~n4045;
  assign n11092 = ~n3805 & n9867;
  assign n11093 = ~n3964 & n10434;
  assign n11094 = ~n11092 & ~n11093;
  assign n11095 = ~n11091 & n11094;
  assign n11096 = n4477 & n9870;
  assign n11097 = n11095 & ~n11096;
  assign n11098 =  a[5]  & ~n11097;
  assign n11099 = ~n11097 & ~n11098;
  assign n11100 =  a[5]  & ~n11098;
  assign n11101 = ~n11099 & ~n11100;
  assign n11102 = ~n11017 & ~n11021;
  assign n11103 = ~n11020 & ~n11021;
  assign n11104 = ~n11102 & ~n11103;
  assign n11105 = ~n11101 & ~n11104;
  assign n11106 = ~n11101 & ~n11105;
  assign n11107 = ~n11104 & ~n11105;
  assign n11108 = ~n11106 & ~n11107;
  assign n11109 = n71 & ~n3964;
  assign n11110 = ~n3456 & n9867;
  assign n11111 = ~n3805 & n10434;
  assign n11112 = ~n11110 & ~n11111;
  assign n11113 = ~n11109 & n11112;
  assign n11114 = n4558 & n9870;
  assign n11115 = n11113 & ~n11114;
  assign n11116 =  a[5]  & ~n11115;
  assign n11117 = ~n11115 & ~n11116;
  assign n11118 =  a[5]  & ~n11116;
  assign n11119 = ~n11117 & ~n11118;
  assign n11120 = ~n11012 & ~n11016;
  assign n11121 = ~n11015 & ~n11016;
  assign n11122 = ~n11120 & ~n11121;
  assign n11123 = ~n11119 & ~n11122;
  assign n11124 = ~n11119 & ~n11123;
  assign n11125 = ~n11122 & ~n11123;
  assign n11126 = ~n11124 & ~n11125;
  assign n11127 = n71 & ~n3805;
  assign n11128 = ~n3605 & n9867;
  assign n11129 = ~n3456 & n10434;
  assign n11130 = ~n11128 & ~n11129;
  assign n11131 = ~n11127 & n11130;
  assign n11132 = n3818 & n9870;
  assign n11133 = n11131 & ~n11132;
  assign n11134 =  a[5]  & ~n11133;
  assign n11135 = ~n11133 & ~n11134;
  assign n11136 =  a[5]  & ~n11134;
  assign n11137 = ~n11135 & ~n11136;
  assign n11138 = ~n11007 & ~n11011;
  assign n11139 = ~n11010 & ~n11011;
  assign n11140 = ~n11138 & ~n11139;
  assign n11141 = ~n11137 & ~n11140;
  assign n11142 = ~n11137 & ~n11141;
  assign n11143 = ~n11140 & ~n11141;
  assign n11144 = ~n11142 & ~n11143;
  assign n11145 = n71 & ~n3456;
  assign n11146 = ~n3539 & n9867;
  assign n11147 = ~n3605 & n10434;
  assign n11148 = ~n11146 & ~n11147;
  assign n11149 = ~n11145 & n11148;
  assign n11150 = n3627 & n9870;
  assign n11151 = n11149 & ~n11150;
  assign n11152 =  a[5]  & ~n11151;
  assign n11153 = ~n11151 & ~n11152;
  assign n11154 =  a[5]  & ~n11152;
  assign n11155 = ~n11153 & ~n11154;
  assign n11156 = ~n11002 & ~n11006;
  assign n11157 = ~n11005 & ~n11006;
  assign n11158 = ~n11156 & ~n11157;
  assign n11159 = ~n11155 & ~n11158;
  assign n11160 = ~n11155 & ~n11159;
  assign n11161 = ~n11158 & ~n11159;
  assign n11162 = ~n11160 & ~n11161;
  assign n11163 = n71 & ~n3605;
  assign n11164 = ~n3012 & n9867;
  assign n11165 = ~n3539 & n10434;
  assign n11166 = ~n11164 & ~n11165;
  assign n11167 = ~n11163 & n11166;
  assign n11168 = n4084 & n9870;
  assign n11169 = n11167 & ~n11168;
  assign n11170 =  a[5]  & ~n11169;
  assign n11171 = ~n11169 & ~n11170;
  assign n11172 =  a[5]  & ~n11170;
  assign n11173 = ~n11171 & ~n11172;
  assign n11174 = ~n10997 & ~n11001;
  assign n11175 = ~n11000 & ~n11001;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = ~n11173 & ~n11176;
  assign n11178 = ~n11173 & ~n11177;
  assign n11179 = ~n11176 & ~n11177;
  assign n11180 = ~n11178 & ~n11179;
  assign n11181 = n71 & ~n3539;
  assign n11182 = ~n392 & n9867;
  assign n11183 = ~n3012 & n10434;
  assign n11184 = ~n11182 & ~n11183;
  assign n11185 = ~n11181 & n11184;
  assign n11186 = n3715 & n9870;
  assign n11187 = n11185 & ~n11186;
  assign n11188 =  a[5]  & ~n11187;
  assign n11189 = ~n11187 & ~n11188;
  assign n11190 =  a[5]  & ~n11188;
  assign n11191 = ~n11189 & ~n11190;
  assign n11192 = ~n10992 & ~n10996;
  assign n11193 = ~n10995 & ~n10996;
  assign n11194 = ~n11192 & ~n11193;
  assign n11195 = ~n11191 & ~n11194;
  assign n11196 = ~n11191 & ~n11195;
  assign n11197 = ~n11194 & ~n11195;
  assign n11198 = ~n11196 & ~n11197;
  assign n11199 = n10568 & n10990;
  assign n11200 = ~n10991 & ~n11199;
  assign n11201 = n71 & ~n3012;
  assign n11202 = ~n587 & n9867;
  assign n11203 = ~n392 & n10434;
  assign n11204 = ~n11202 & ~n11203;
  assign n11205 = ~n11201 & n11204;
  assign n11206 = ~n9870 & n11205;
  assign n11207 = ~n3018 & n11205;
  assign n11208 = ~n11206 & ~n11207;
  assign n11209 =  a[5]  & ~n11208;
  assign n11210 = ~ a[5]  & n11208;
  assign n11211 = ~n11209 & ~n11210;
  assign n11212 = n11200 & ~n11211;
  assign n11213 = n10586 & n10988;
  assign n11214 = ~n10989 & ~n11213;
  assign n11215 = n71 & ~n392;
  assign n11216 = ~n710 & n9867;
  assign n11217 = ~n587 & n10434;
  assign n11218 = ~n11216 & ~n11217;
  assign n11219 = ~n11215 & n11218;
  assign n11220 = ~n9870 & n11219;
  assign n11221 = ~n3347 & n11219;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 =  a[5]  & ~n11222;
  assign n11224 = ~ a[5]  & n11222;
  assign n11225 = ~n11223 & ~n11224;
  assign n11226 = n11214 & ~n11225;
  assign n11227 = n71 & ~n587;
  assign n11228 = ~n867 & n9867;
  assign n11229 = ~n710 & n10434;
  assign n11230 = ~n11228 & ~n11229;
  assign n11231 = ~n11227 & n11230;
  assign n11232 = n3331 & n9870;
  assign n11233 = n11231 & ~n11232;
  assign n11234 =  a[5]  & ~n11233;
  assign n11235 = ~n11233 & ~n11234;
  assign n11236 =  a[5]  & ~n11234;
  assign n11237 = ~n11235 & ~n11236;
  assign n11238 = n10984 & ~n10986;
  assign n11239 = ~n10987 & ~n11238;
  assign n11240 = ~n11237 & n11239;
  assign n11241 = ~n11237 & ~n11240;
  assign n11242 = n11239 & ~n11240;
  assign n11243 = ~n11241 & ~n11242;
  assign n11244 = n71 & ~n710;
  assign n11245 = ~n958 & n9867;
  assign n11246 = ~n867 & n10434;
  assign n11247 = ~n11245 & ~n11246;
  assign n11248 = ~n11244 & n11247;
  assign n11249 = n4179 & n9870;
  assign n11250 = n11248 & ~n11249;
  assign n11251 =  a[5]  & ~n11250;
  assign n11252 = ~n11250 & ~n11251;
  assign n11253 =  a[5]  & ~n11251;
  assign n11254 = ~n11252 & ~n11253;
  assign n11255 = ~n10979 & ~n10983;
  assign n11256 = ~n10982 & ~n10983;
  assign n11257 = ~n11255 & ~n11256;
  assign n11258 = ~n11254 & ~n11257;
  assign n11259 = ~n11254 & ~n11258;
  assign n11260 = ~n11257 & ~n11258;
  assign n11261 = ~n11259 & ~n11260;
  assign n11262 = n71 & ~n867;
  assign n11263 = ~n1060 & n9867;
  assign n11264 = ~n958 & n10434;
  assign n11265 = ~n11263 & ~n11264;
  assign n11266 = ~n11262 & n11265;
  assign n11267 = n4204 & n9870;
  assign n11268 = n11266 & ~n11267;
  assign n11269 =  a[5]  & ~n11268;
  assign n11270 = ~n11268 & ~n11269;
  assign n11271 =  a[5]  & ~n11269;
  assign n11272 = ~n11270 & ~n11271;
  assign n11273 = ~n10974 & ~n10978;
  assign n11274 = ~n10977 & ~n10978;
  assign n11275 = ~n11273 & ~n11274;
  assign n11276 = ~n11272 & ~n11275;
  assign n11277 = ~n11272 & ~n11276;
  assign n11278 = ~n11275 & ~n11276;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = n10645 & n10972;
  assign n11281 = ~n10973 & ~n11280;
  assign n11282 = n71 & ~n958;
  assign n11283 = ~n1178 & n9867;
  assign n11284 = ~n1060 & n10434;
  assign n11285 = ~n11283 & ~n11284;
  assign n11286 = ~n11282 & n11285;
  assign n11287 = ~n9870 & n11286;
  assign n11288 = ~n4633 & n11286;
  assign n11289 = ~n11287 & ~n11288;
  assign n11290 =  a[5]  & ~n11289;
  assign n11291 = ~ a[5]  & n11289;
  assign n11292 = ~n11290 & ~n11291;
  assign n11293 = n11281 & ~n11292;
  assign n11294 = n10663 & n10970;
  assign n11295 = ~n10971 & ~n11294;
  assign n11296 = n71 & ~n1060;
  assign n11297 = ~n1235 & n9867;
  assign n11298 = ~n1178 & n10434;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = ~n11296 & n11299;
  assign n11301 = ~n9870 & n11300;
  assign n11302 = ~n4429 & n11300;
  assign n11303 = ~n11301 & ~n11302;
  assign n11304 =  a[5]  & ~n11303;
  assign n11305 = ~ a[5]  & n11303;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = n11295 & ~n11306;
  assign n11308 = n10681 & n10968;
  assign n11309 = ~n10969 & ~n11308;
  assign n11310 = n71 & ~n1178;
  assign n11311 = ~n1364 & n9867;
  assign n11312 = ~n1235 & n10434;
  assign n11313 = ~n11311 & ~n11312;
  assign n11314 = ~n11310 & n11313;
  assign n11315 = ~n9870 & n11314;
  assign n11316 = ~n4861 & n11314;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 =  a[5]  & ~n11317;
  assign n11319 = ~ a[5]  & n11317;
  assign n11320 = ~n11318 & ~n11319;
  assign n11321 = n11309 & ~n11320;
  assign n11322 = n71 & ~n1235;
  assign n11323 = ~n1472 & n9867;
  assign n11324 = ~n1364 & n10434;
  assign n11325 = ~n11323 & ~n11324;
  assign n11326 = ~n11322 & n11325;
  assign n11327 = n4848 & n9870;
  assign n11328 = n11326 & ~n11327;
  assign n11329 =  a[5]  & ~n11328;
  assign n11330 = ~n11328 & ~n11329;
  assign n11331 =  a[5]  & ~n11329;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = n10964 & ~n10966;
  assign n11334 = ~n10967 & ~n11333;
  assign n11335 = ~n11332 & n11334;
  assign n11336 = ~n11332 & ~n11335;
  assign n11337 = n11334 & ~n11335;
  assign n11338 = ~n11336 & ~n11337;
  assign n11339 = n71 & ~n1364;
  assign n11340 = ~n1572 & n9867;
  assign n11341 = ~n1472 & n10434;
  assign n11342 = ~n11340 & ~n11341;
  assign n11343 = ~n11339 & n11342;
  assign n11344 = n5114 & n9870;
  assign n11345 = n11343 & ~n11344;
  assign n11346 =  a[5]  & ~n11345;
  assign n11347 = ~n11345 & ~n11346;
  assign n11348 =  a[5]  & ~n11346;
  assign n11349 = ~n11347 & ~n11348;
  assign n11350 = ~n10959 & ~n10963;
  assign n11351 = ~n10962 & ~n10963;
  assign n11352 = ~n11350 & ~n11351;
  assign n11353 = ~n11349 & ~n11352;
  assign n11354 = ~n11349 & ~n11353;
  assign n11355 = ~n11352 & ~n11353;
  assign n11356 = ~n11354 & ~n11355;
  assign n11357 = n71 & ~n1472;
  assign n11358 = ~n1665 & n9867;
  assign n11359 = ~n1572 & n10434;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = ~n11357 & n11360;
  assign n11362 = n5139 & n9870;
  assign n11363 = n11361 & ~n11362;
  assign n11364 =  a[5]  & ~n11363;
  assign n11365 = ~n11363 & ~n11364;
  assign n11366 =  a[5]  & ~n11364;
  assign n11367 = ~n11365 & ~n11366;
  assign n11368 = ~n10954 & ~n10958;
  assign n11369 = ~n10957 & ~n10958;
  assign n11370 = ~n11368 & ~n11369;
  assign n11371 = ~n11367 & ~n11370;
  assign n11372 = ~n11367 & ~n11371;
  assign n11373 = ~n11370 & ~n11371;
  assign n11374 = ~n11372 & ~n11373;
  assign n11375 = n10740 & n10952;
  assign n11376 = ~n10953 & ~n11375;
  assign n11377 = n71 & ~n1572;
  assign n11378 = ~n1779 & n9867;
  assign n11379 = ~n1665 & n10434;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = ~n11377 & n11380;
  assign n11382 = ~n9870 & n11381;
  assign n11383 = ~n5561 & n11381;
  assign n11384 = ~n11382 & ~n11383;
  assign n11385 =  a[5]  & ~n11384;
  assign n11386 = ~ a[5]  & n11384;
  assign n11387 = ~n11385 & ~n11386;
  assign n11388 = n11376 & ~n11387;
  assign n11389 = n10758 & n10950;
  assign n11390 = ~n10951 & ~n11389;
  assign n11391 = n71 & ~n1665;
  assign n11392 = ~n1877 & n9867;
  assign n11393 = ~n1779 & n10434;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = ~n11391 & n11394;
  assign n11396 = ~n9870 & n11395;
  assign n11397 = ~n5328 & n11395;
  assign n11398 = ~n11396 & ~n11397;
  assign n11399 =  a[5]  & ~n11398;
  assign n11400 = ~ a[5]  & n11398;
  assign n11401 = ~n11399 & ~n11400;
  assign n11402 = n11390 & ~n11401;
  assign n11403 = n10776 & n10948;
  assign n11404 = ~n10949 & ~n11403;
  assign n11405 = n71 & ~n1779;
  assign n11406 = ~n1913 & n9867;
  assign n11407 = ~n1877 & n10434;
  assign n11408 = ~n11406 & ~n11407;
  assign n11409 = ~n11405 & n11408;
  assign n11410 = ~n9870 & n11409;
  assign n11411 = ~n5851 & n11409;
  assign n11412 = ~n11410 & ~n11411;
  assign n11413 =  a[5]  & ~n11412;
  assign n11414 = ~ a[5]  & n11412;
  assign n11415 = ~n11413 & ~n11414;
  assign n11416 = n11404 & ~n11415;
  assign n11417 = n71 & ~n1877;
  assign n11418 = ~n1992 & n9867;
  assign n11419 = ~n1913 & n10434;
  assign n11420 = ~n11418 & ~n11419;
  assign n11421 = ~n11417 & n11420;
  assign n11422 = n6007 & n9870;
  assign n11423 = n11421 & ~n11422;
  assign n11424 =  a[5]  & ~n11423;
  assign n11425 = ~n11423 & ~n11424;
  assign n11426 =  a[5]  & ~n11424;
  assign n11427 = ~n11425 & ~n11426;
  assign n11428 = n10944 & ~n10946;
  assign n11429 = ~n10947 & ~n11428;
  assign n11430 = ~n11427 & n11429;
  assign n11431 = ~n11427 & ~n11430;
  assign n11432 = n11429 & ~n11430;
  assign n11433 = ~n11431 & ~n11432;
  assign n11434 = n71 & ~n1913;
  assign n11435 = ~n2057 & n9867;
  assign n11436 = ~n1992 & n10434;
  assign n11437 = ~n11435 & ~n11436;
  assign n11438 = ~n11434 & n11437;
  assign n11439 = n5834 & n9870;
  assign n11440 = n11438 & ~n11439;
  assign n11441 =  a[5]  & ~n11440;
  assign n11442 = ~n11440 & ~n11441;
  assign n11443 =  a[5]  & ~n11441;
  assign n11444 = ~n11442 & ~n11443;
  assign n11445 = ~n10939 & ~n10943;
  assign n11446 = ~n10942 & ~n10943;
  assign n11447 = ~n11445 & ~n11446;
  assign n11448 = ~n11444 & ~n11447;
  assign n11449 = ~n11444 & ~n11448;
  assign n11450 = ~n11447 & ~n11448;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = n71 & ~n1992;
  assign n11453 = ~n2152 & n9867;
  assign n11454 = ~n2057 & n10434;
  assign n11455 = ~n11453 & ~n11454;
  assign n11456 = ~n11452 & n11455;
  assign n11457 = n6143 & n9870;
  assign n11458 = n11456 & ~n11457;
  assign n11459 =  a[5]  & ~n11458;
  assign n11460 = ~n11458 & ~n11459;
  assign n11461 =  a[5]  & ~n11459;
  assign n11462 = ~n11460 & ~n11461;
  assign n11463 = ~n10934 & ~n10938;
  assign n11464 = ~n10937 & ~n10938;
  assign n11465 = ~n11463 & ~n11464;
  assign n11466 = ~n11462 & ~n11465;
  assign n11467 = ~n11462 & ~n11466;
  assign n11468 = ~n11465 & ~n11466;
  assign n11469 = ~n11467 & ~n11468;
  assign n11470 = n10835 & n10932;
  assign n11471 = ~n10933 & ~n11470;
  assign n11472 = n71 & ~n2057;
  assign n11473 = ~n2189 & n9867;
  assign n11474 = ~n2152 & n10434;
  assign n11475 = ~n11473 & ~n11474;
  assign n11476 = ~n11472 & n11475;
  assign n11477 = ~n9870 & n11476;
  assign n11478 = ~n6479 & n11476;
  assign n11479 = ~n11477 & ~n11478;
  assign n11480 =  a[5]  & ~n11479;
  assign n11481 = ~ a[5]  & n11479;
  assign n11482 = ~n11480 & ~n11481;
  assign n11483 = n11471 & ~n11482;
  assign n11484 = n10928 & ~n10930;
  assign n11485 = ~n10931 & ~n11484;
  assign n11486 = n71 & ~n2152;
  assign n11487 = ~n2291 & n9867;
  assign n11488 = ~n2189 & n10434;
  assign n11489 = ~n11487 & ~n11488;
  assign n11490 = ~n11486 & n11489;
  assign n11491 = ~n9870 & n11490;
  assign n11492 = ~n6492 & n11490;
  assign n11493 = ~n11491 & ~n11492;
  assign n11494 =  a[5]  & ~n11493;
  assign n11495 = ~ a[5]  & n11493;
  assign n11496 = ~n11494 & ~n11495;
  assign n11497 = n11485 & ~n11496;
  assign n11498 = n10867 & n10926;
  assign n11499 = ~n10927 & ~n11498;
  assign n11500 = n71 & ~n2189;
  assign n11501 = ~n2388 & n9867;
  assign n11502 = ~n2291 & n10434;
  assign n11503 = ~n11501 & ~n11502;
  assign n11504 = ~n11500 & n11503;
  assign n11505 = ~n9870 & n11504;
  assign n11506 = ~n6122 & n11504;
  assign n11507 = ~n11505 & ~n11506;
  assign n11508 =  a[5]  & ~n11507;
  assign n11509 = ~ a[5]  & n11507;
  assign n11510 = ~n11508 & ~n11509;
  assign n11511 = n11499 & ~n11510;
  assign n11512 = n71 & ~n2291;
  assign n11513 = ~n2464 & n9867;
  assign n11514 = ~n2388 & n10434;
  assign n11515 = ~n11513 & ~n11514;
  assign n11516 = ~n11512 & n11515;
  assign n11517 = n6541 & n9870;
  assign n11518 = n11516 & ~n11517;
  assign n11519 =  a[5]  & ~n11518;
  assign n11520 = ~n11518 & ~n11519;
  assign n11521 =  a[5]  & ~n11519;
  assign n11522 = ~n11520 & ~n11521;
  assign n11523 = n10922 & ~n10924;
  assign n11524 = ~n10925 & ~n11523;
  assign n11525 = ~n11522 & n11524;
  assign n11526 = ~n11522 & ~n11525;
  assign n11527 = n11524 & ~n11525;
  assign n11528 = ~n11526 & ~n11527;
  assign n11529 = ~n10909 & ~n10921;
  assign n11530 = ~n10920 & ~n10921;
  assign n11531 = ~n11529 & ~n11530;
  assign n11532 = n71 & ~n2388;
  assign n11533 = ~n2533 & n9867;
  assign n11534 = ~n2464 & n10434;
  assign n11535 = ~n11533 & ~n11534;
  assign n11536 = ~n11532 & n11535;
  assign n11537 = ~n9870 & n11536;
  assign n11538 = ~n6591 & n11536;
  assign n11539 = ~n11537 & ~n11538;
  assign n11540 =  a[5]  & ~n11539;
  assign n11541 = ~ a[5]  & n11539;
  assign n11542 = ~n11540 & ~n11541;
  assign n11543 = ~n11531 & ~n11542;
  assign n11544 = n71 & ~n2464;
  assign n11545 = ~n2571 & n9867;
  assign n11546 = ~n2533 & n10434;
  assign n11547 = ~n11545 & ~n11546;
  assign n11548 = ~n11544 & n11547;
  assign n11549 = n6646 & n9870;
  assign n11550 = n11548 & ~n11549;
  assign n11551 =  a[5]  & ~n11550;
  assign n11552 = ~n11550 & ~n11551;
  assign n11553 =  a[5]  & ~n11551;
  assign n11554 = ~n11552 & ~n11553;
  assign n11555 = ~n10893 & n10904;
  assign n11556 = ~n10905 & ~n11555;
  assign n11557 = ~n11554 & n11556;
  assign n11558 = ~n11554 & ~n11557;
  assign n11559 = n11556 & ~n11557;
  assign n11560 = ~n11558 & ~n11559;
  assign n11561 = n10890 & ~n10892;
  assign n11562 = ~n10893 & ~n11561;
  assign n11563 = n71 & ~n2533;
  assign n11564 = ~n2674 & n9867;
  assign n11565 = ~n2571 & n10434;
  assign n11566 = ~n11564 & ~n11565;
  assign n11567 = ~n11563 & n11566;
  assign n11568 = ~n9870 & n11567;
  assign n11569 = ~n6695 & n11567;
  assign n11570 = ~n11568 & ~n11569;
  assign n11571 =  a[5]  & ~n11570;
  assign n11572 = ~ a[5]  & n11570;
  assign n11573 = ~n11571 & ~n11572;
  assign n11574 = n11562 & ~n11573;
  assign n11575 = ~n2829 & n10434;
  assign n11576 = n71 & ~n2736;
  assign n11577 = ~n11575 & ~n11576;
  assign n11578 = ~n7469 & n9870;
  assign n11579 = n11577 & ~n11578;
  assign n11580 =  a[5]  & ~n11579;
  assign n11581 =  a[5]  & ~n11580;
  assign n11582 = ~n11579 & ~n11580;
  assign n11583 = ~n11581 & ~n11582;
  assign n11584 = ~n70 & ~n2829;
  assign n11585 =  a[5]  & ~n11584;
  assign n11586 = ~n11583 & n11585;
  assign n11587 = n71 & ~n2674;
  assign n11588 = ~n2829 & n9867;
  assign n11589 = ~n2736 & n10434;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = ~n11587 & n11590;
  assign n11592 = ~n9870 & n11591;
  assign n11593 = ~n6798 & n11591;
  assign n11594 = ~n11592 & ~n11593;
  assign n11595 =  a[5]  & ~n11594;
  assign n11596 = ~ a[5]  & n11594;
  assign n11597 = ~n11595 & ~n11596;
  assign n11598 = n11586 & ~n11597;
  assign n11599 = n10891 & n11598;
  assign n11600 = n11598 & ~n11599;
  assign n11601 = n10891 & ~n11599;
  assign n11602 = ~n11600 & ~n11601;
  assign n11603 = n71 & ~n2571;
  assign n11604 = ~n2736 & n9867;
  assign n11605 = ~n2674 & n10434;
  assign n11606 = ~n11604 & ~n11605;
  assign n11607 = ~n11603 & n11606;
  assign n11608 = n6806 & n9870;
  assign n11609 = n11607 & ~n11608;
  assign n11610 =  a[5]  & ~n11609;
  assign n11611 =  a[5]  & ~n11610;
  assign n11612 = ~n11609 & ~n11610;
  assign n11613 = ~n11611 & ~n11612;
  assign n11614 = ~n11602 & ~n11613;
  assign n11615 = ~n11599 & ~n11614;
  assign n11616 = ~n11562 & n11573;
  assign n11617 = ~n11574 & ~n11616;
  assign n11618 = ~n11615 & n11617;
  assign n11619 = ~n11574 & ~n11618;
  assign n11620 = ~n11560 & ~n11619;
  assign n11621 = ~n11557 & ~n11620;
  assign n11622 = n11531 & n11542;
  assign n11623 = ~n11543 & ~n11622;
  assign n11624 = ~n11621 & n11623;
  assign n11625 = ~n11543 & ~n11624;
  assign n11626 = ~n11528 & ~n11625;
  assign n11627 = ~n11525 & ~n11626;
  assign n11628 = n11499 & ~n11511;
  assign n11629 = ~n11510 & ~n11511;
  assign n11630 = ~n11628 & ~n11629;
  assign n11631 = ~n11627 & ~n11630;
  assign n11632 = ~n11511 & ~n11631;
  assign n11633 = n11485 & ~n11497;
  assign n11634 = ~n11496 & ~n11497;
  assign n11635 = ~n11633 & ~n11634;
  assign n11636 = ~n11632 & ~n11635;
  assign n11637 = ~n11497 & ~n11636;
  assign n11638 = ~n11471 & n11482;
  assign n11639 = ~n11483 & ~n11638;
  assign n11640 = ~n11637 & n11639;
  assign n11641 = ~n11483 & ~n11640;
  assign n11642 = ~n11469 & ~n11641;
  assign n11643 = ~n11466 & ~n11642;
  assign n11644 = ~n11451 & ~n11643;
  assign n11645 = ~n11448 & ~n11644;
  assign n11646 = ~n11433 & ~n11645;
  assign n11647 = ~n11430 & ~n11646;
  assign n11648 = n11404 & ~n11416;
  assign n11649 = ~n11415 & ~n11416;
  assign n11650 = ~n11648 & ~n11649;
  assign n11651 = ~n11647 & ~n11650;
  assign n11652 = ~n11416 & ~n11651;
  assign n11653 = n11390 & ~n11402;
  assign n11654 = ~n11401 & ~n11402;
  assign n11655 = ~n11653 & ~n11654;
  assign n11656 = ~n11652 & ~n11655;
  assign n11657 = ~n11402 & ~n11656;
  assign n11658 = ~n11376 & n11387;
  assign n11659 = ~n11388 & ~n11658;
  assign n11660 = ~n11657 & n11659;
  assign n11661 = ~n11388 & ~n11660;
  assign n11662 = ~n11374 & ~n11661;
  assign n11663 = ~n11371 & ~n11662;
  assign n11664 = ~n11356 & ~n11663;
  assign n11665 = ~n11353 & ~n11664;
  assign n11666 = ~n11338 & ~n11665;
  assign n11667 = ~n11335 & ~n11666;
  assign n11668 = n11309 & ~n11321;
  assign n11669 = ~n11320 & ~n11321;
  assign n11670 = ~n11668 & ~n11669;
  assign n11671 = ~n11667 & ~n11670;
  assign n11672 = ~n11321 & ~n11671;
  assign n11673 = n11295 & ~n11307;
  assign n11674 = ~n11306 & ~n11307;
  assign n11675 = ~n11673 & ~n11674;
  assign n11676 = ~n11672 & ~n11675;
  assign n11677 = ~n11307 & ~n11676;
  assign n11678 = ~n11281 & n11292;
  assign n11679 = ~n11293 & ~n11678;
  assign n11680 = ~n11677 & n11679;
  assign n11681 = ~n11293 & ~n11680;
  assign n11682 = ~n11279 & ~n11681;
  assign n11683 = ~n11276 & ~n11682;
  assign n11684 = ~n11261 & ~n11683;
  assign n11685 = ~n11258 & ~n11684;
  assign n11686 = ~n11243 & ~n11685;
  assign n11687 = ~n11240 & ~n11686;
  assign n11688 = n11214 & ~n11226;
  assign n11689 = ~n11225 & ~n11226;
  assign n11690 = ~n11688 & ~n11689;
  assign n11691 = ~n11687 & ~n11690;
  assign n11692 = ~n11226 & ~n11691;
  assign n11693 = ~n11200 & n11211;
  assign n11694 = ~n11212 & ~n11693;
  assign n11695 = ~n11692 & n11694;
  assign n11696 = ~n11212 & ~n11695;
  assign n11697 = ~n11198 & ~n11696;
  assign n11698 = ~n11195 & ~n11697;
  assign n11699 = ~n11180 & ~n11698;
  assign n11700 = ~n11177 & ~n11699;
  assign n11701 = ~n11162 & ~n11700;
  assign n11702 = ~n11159 & ~n11701;
  assign n11703 = ~n11144 & ~n11702;
  assign n11704 = ~n11141 & ~n11703;
  assign n11705 = ~n11126 & ~n11704;
  assign n11706 = ~n11123 & ~n11705;
  assign n11707 = ~n11108 & ~n11706;
  assign n11708 = ~n11105 & ~n11707;
  assign n11709 = ~n11090 & ~n11708;
  assign n11710 = n11090 & n11708;
  assign n11711 = ~n11709 & ~n11710;
  assign n11712 = n11108 & n11706;
  assign n11713 = ~n11707 & ~n11712;
  assign n11714 = ~n3877 & n11055;
  assign n11715 = ~ a[0]  &  a[1] ;
  assign n11716 = ~n4515 & n11715;
  assign n11717 = ~n11714 & ~n11716;
  assign n11718 = ~n11057 & n11717;
  assign n11719 = ~n4609 & n11717;
  assign n11720 = ~n11718 & ~n11719;
  assign n11721 =  a[2]  & ~n11720;
  assign n11722 = ~ a[2]  & n11720;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = n11713 & ~n11723;
  assign n11725 = n11126 & n11704;
  assign n11726 = ~n11705 & ~n11725;
  assign n11727 =  a[0]  & n11053;
  assign n11728 = ~n4515 & n11727;
  assign n11729 = ~n4045 & n11055;
  assign n11730 = ~n3877 & n11715;
  assign n11731 = ~n11729 & ~n11730;
  assign n11732 = ~n11728 & n11731;
  assign n11733 = ~n11057 & n11732;
  assign n11734 = ~n4715 & n11732;
  assign n11735 = ~n11733 & ~n11734;
  assign n11736 =  a[2]  & ~n11735;
  assign n11737 = ~ a[2]  & n11735;
  assign n11738 = ~n11736 & ~n11737;
  assign n11739 = n11726 & ~n11738;
  assign n11740 = n11144 & n11702;
  assign n11741 = ~n11703 & ~n11740;
  assign n11742 = ~n3877 & n11727;
  assign n11743 = ~n3964 & n11055;
  assign n11744 = ~n4045 & n11715;
  assign n11745 = ~n11743 & ~n11744;
  assign n11746 = ~n11742 & n11745;
  assign n11747 = ~n11057 & n11746;
  assign n11748 = ~n4067 & n11746;
  assign n11749 = ~n11747 & ~n11748;
  assign n11750 =  a[2]  & ~n11749;
  assign n11751 = ~ a[2]  & n11749;
  assign n11752 = ~n11750 & ~n11751;
  assign n11753 = n11741 & ~n11752;
  assign n11754 = n11162 & n11700;
  assign n11755 = ~n11701 & ~n11754;
  assign n11756 = ~n4045 & n11727;
  assign n11757 = ~n3805 & n11055;
  assign n11758 = ~n3964 & n11715;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = ~n11756 & n11759;
  assign n11761 = ~n11057 & n11760;
  assign n11762 = ~n4477 & n11760;
  assign n11763 = ~n11761 & ~n11762;
  assign n11764 =  a[2]  & ~n11763;
  assign n11765 = ~ a[2]  & n11763;
  assign n11766 = ~n11764 & ~n11765;
  assign n11767 = n11755 & ~n11766;
  assign n11768 = n11180 & n11698;
  assign n11769 = ~n11699 & ~n11768;
  assign n11770 = ~n3964 & n11727;
  assign n11771 = ~n3456 & n11055;
  assign n11772 = ~n3805 & n11715;
  assign n11773 = ~n11771 & ~n11772;
  assign n11774 = ~n11770 & n11773;
  assign n11775 = ~n11057 & n11774;
  assign n11776 = ~n4558 & n11774;
  assign n11777 = ~n11775 & ~n11776;
  assign n11778 =  a[2]  & ~n11777;
  assign n11779 = ~ a[2]  & n11777;
  assign n11780 = ~n11778 & ~n11779;
  assign n11781 = n11769 & ~n11780;
  assign n11782 = n11692 & ~n11694;
  assign n11783 = ~n11695 & ~n11782;
  assign n11784 = n11677 & ~n11679;
  assign n11785 = ~n11680 & ~n11784;
  assign n11786 = n11657 & ~n11659;
  assign n11787 = ~n11660 & ~n11786;
  assign n11788 = n11637 & ~n11639;
  assign n11789 = ~n11640 & ~n11788;
  assign n11790 = n11615 & ~n11617;
  assign n11791 = ~n11618 & ~n11790;
  assign n11792 = ~n11586 & n11597;
  assign n11793 = ~n11598 & ~n11792;
  assign n11794 = ~n11057 & ~n11727;
  assign n11795 = ~n2829 & ~n11794;
  assign n11796 =  a[2]  & n11057;
  assign n11797 = n6798 & n11796;
  assign n11798 = ~n2674 & n11727;
  assign n11799 = ~n2829 & n11055;
  assign n11800 = ~n2736 & n11715;
  assign n11801 = ~n11799 & ~n11800;
  assign n11802 = ~n11798 & n11801;
  assign n11803 =  a[2]  & ~n11802;
  assign n11804 = ~n7469 & n11796;
  assign n11805 =  a[2]  & n11715;
  assign n11806 = ~n2829 & n11805;
  assign n11807 =  a[2]  & n11727;
  assign n11808 = ~n2736 & n11807;
  assign n11809 =  a[2]  & ~n11808;
  assign n11810 = ~n11806 & n11809;
  assign n11811 = ~n11804 & n11810;
  assign n11812 = ~n11803 & n11811;
  assign n11813 = ~n11797 & n11812;
  assign n11814 = ~n11795 & n11813;
  assign n11815 = n11584 & n11814;
  assign n11816 = ~n11584 & ~n11814;
  assign n11817 = ~n2571 & n11727;
  assign n11818 = ~n2736 & n11055;
  assign n11819 = ~n2674 & n11715;
  assign n11820 = ~n11818 & ~n11819;
  assign n11821 = ~n11817 & n11820;
  assign n11822 = n6806 & n11057;
  assign n11823 = n11821 & ~n11822;
  assign n11824 = ~ a[2]  & ~n11823;
  assign n11825 =  a[2]  & n11823;
  assign n11826 = ~n11824 & ~n11825;
  assign n11827 = ~n11816 & ~n11826;
  assign n11828 = ~n11815 & ~n11827;
  assign n11829 = ~n2533 & n11727;
  assign n11830 = ~n2674 & n11055;
  assign n11831 = ~n2571 & n11715;
  assign n11832 = ~n11830 & ~n11831;
  assign n11833 = ~n11829 & n11832;
  assign n11834 = ~n11057 & n11833;
  assign n11835 = ~n6695 & n11833;
  assign n11836 = ~n11834 & ~n11835;
  assign n11837 =  a[2]  & ~n11836;
  assign n11838 = ~ a[2]  & n11836;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = n11828 & n11839;
  assign n11841 = n11583 & ~n11585;
  assign n11842 = ~n11586 & ~n11841;
  assign n11843 = ~n11840 & n11842;
  assign n11844 = ~n11828 & ~n11839;
  assign n11845 = ~n11843 & ~n11844;
  assign n11846 = n11793 & ~n11845;
  assign n11847 = ~n11793 & n11845;
  assign n11848 = ~n2464 & n11727;
  assign n11849 = ~n2571 & n11055;
  assign n11850 = ~n2533 & n11715;
  assign n11851 = ~n11849 & ~n11850;
  assign n11852 = ~n11848 & n11851;
  assign n11853 = n6646 & n11057;
  assign n11854 = n11852 & ~n11853;
  assign n11855 = ~ a[2]  & ~n11854;
  assign n11856 =  a[2]  & n11854;
  assign n11857 = ~n11855 & ~n11856;
  assign n11858 = ~n11847 & ~n11857;
  assign n11859 = ~n11846 & ~n11858;
  assign n11860 = ~n2388 & n11727;
  assign n11861 = ~n2533 & n11055;
  assign n11862 = ~n2464 & n11715;
  assign n11863 = ~n11861 & ~n11862;
  assign n11864 = ~n11860 & n11863;
  assign n11865 = ~n11057 & n11864;
  assign n11866 = ~n6591 & n11864;
  assign n11867 = ~n11865 & ~n11866;
  assign n11868 =  a[2]  & ~n11867;
  assign n11869 = ~ a[2]  & n11867;
  assign n11870 = ~n11868 & ~n11869;
  assign n11871 = ~n11859 & ~n11870;
  assign n11872 = n11859 & n11870;
  assign n11873 = n11602 & n11613;
  assign n11874 = ~n11614 & ~n11873;
  assign n11875 = ~n11872 & n11874;
  assign n11876 = ~n11871 & ~n11875;
  assign n11877 = n11791 & ~n11876;
  assign n11878 = ~n11791 & n11876;
  assign n11879 = ~n2291 & n11727;
  assign n11880 = ~n2464 & n11055;
  assign n11881 = ~n2388 & n11715;
  assign n11882 = ~n11880 & ~n11881;
  assign n11883 = ~n11879 & n11882;
  assign n11884 = n6541 & n11057;
  assign n11885 = n11883 & ~n11884;
  assign n11886 = ~ a[2]  & ~n11885;
  assign n11887 =  a[2]  & n11885;
  assign n11888 = ~n11886 & ~n11887;
  assign n11889 = ~n11878 & ~n11888;
  assign n11890 = ~n11877 & ~n11889;
  assign n11891 = ~n2189 & n11727;
  assign n11892 = ~n2388 & n11055;
  assign n11893 = ~n2291 & n11715;
  assign n11894 = ~n11892 & ~n11893;
  assign n11895 = ~n11891 & n11894;
  assign n11896 = ~n11057 & n11895;
  assign n11897 = ~n6122 & n11895;
  assign n11898 = ~n11896 & ~n11897;
  assign n11899 =  a[2]  & ~n11898;
  assign n11900 = ~ a[2]  & n11898;
  assign n11901 = ~n11899 & ~n11900;
  assign n11902 = n11890 & n11901;
  assign n11903 = n11560 & n11619;
  assign n11904 = ~n11620 & ~n11903;
  assign n11905 = ~n11902 & n11904;
  assign n11906 = ~n11890 & ~n11901;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = ~n2152 & n11727;
  assign n11909 = ~n2291 & n11055;
  assign n11910 = ~n2189 & n11715;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = ~n11908 & n11911;
  assign n11913 = ~n11057 & n11912;
  assign n11914 = ~n6492 & n11912;
  assign n11915 = ~n11913 & ~n11914;
  assign n11916 =  a[2]  & ~n11915;
  assign n11917 = ~ a[2]  & n11915;
  assign n11918 = ~n11916 & ~n11917;
  assign n11919 = n11907 & n11918;
  assign n11920 = n11621 & ~n11623;
  assign n11921 = ~n11624 & ~n11920;
  assign n11922 = ~n11919 & n11921;
  assign n11923 = ~n11907 & ~n11918;
  assign n11924 = ~n11922 & ~n11923;
  assign n11925 = ~n2057 & n11727;
  assign n11926 = ~n2189 & n11055;
  assign n11927 = ~n2152 & n11715;
  assign n11928 = ~n11926 & ~n11927;
  assign n11929 = ~n11925 & n11928;
  assign n11930 = ~n11057 & n11929;
  assign n11931 = ~n6479 & n11929;
  assign n11932 = ~n11930 & ~n11931;
  assign n11933 =  a[2]  & ~n11932;
  assign n11934 = ~ a[2]  & n11932;
  assign n11935 = ~n11933 & ~n11934;
  assign n11936 = n11924 & n11935;
  assign n11937 = n11528 & n11625;
  assign n11938 = ~n11626 & ~n11937;
  assign n11939 = ~n11936 & n11938;
  assign n11940 = ~n11924 & ~n11935;
  assign n11941 = ~n11939 & ~n11940;
  assign n11942 = n11627 & ~n11629;
  assign n11943 = ~n11628 & n11942;
  assign n11944 = ~n11631 & ~n11943;
  assign n11945 = ~n11941 & n11944;
  assign n11946 = n11941 & ~n11944;
  assign n11947 = ~n1992 & n11727;
  assign n11948 = ~n2152 & n11055;
  assign n11949 = ~n2057 & n11715;
  assign n11950 = ~n11948 & ~n11949;
  assign n11951 = ~n11947 & n11950;
  assign n11952 = n6143 & n11057;
  assign n11953 = n11951 & ~n11952;
  assign n11954 = ~ a[2]  & ~n11953;
  assign n11955 =  a[2]  & n11953;
  assign n11956 = ~n11954 & ~n11955;
  assign n11957 = ~n11946 & ~n11956;
  assign n11958 = ~n11945 & ~n11957;
  assign n11959 = n11632 & ~n11634;
  assign n11960 = ~n11633 & n11959;
  assign n11961 = ~n11636 & ~n11960;
  assign n11962 = ~n11958 & n11961;
  assign n11963 = n11958 & ~n11961;
  assign n11964 = ~n1913 & n11727;
  assign n11965 = ~n2057 & n11055;
  assign n11966 = ~n1992 & n11715;
  assign n11967 = ~n11965 & ~n11966;
  assign n11968 = ~n11964 & n11967;
  assign n11969 = n5834 & n11057;
  assign n11970 = n11968 & ~n11969;
  assign n11971 = ~ a[2]  & ~n11970;
  assign n11972 =  a[2]  & n11970;
  assign n11973 = ~n11971 & ~n11972;
  assign n11974 = ~n11963 & ~n11973;
  assign n11975 = ~n11962 & ~n11974;
  assign n11976 = n11789 & ~n11975;
  assign n11977 = ~n11789 & n11975;
  assign n11978 = ~n1877 & n11727;
  assign n11979 = ~n1992 & n11055;
  assign n11980 = ~n1913 & n11715;
  assign n11981 = ~n11979 & ~n11980;
  assign n11982 = ~n11978 & n11981;
  assign n11983 = n6007 & n11057;
  assign n11984 = n11982 & ~n11983;
  assign n11985 = ~ a[2]  & ~n11984;
  assign n11986 =  a[2]  & n11984;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = ~n11977 & ~n11987;
  assign n11989 = ~n11976 & ~n11988;
  assign n11990 = ~n1779 & n11727;
  assign n11991 = ~n1913 & n11055;
  assign n11992 = ~n1877 & n11715;
  assign n11993 = ~n11991 & ~n11992;
  assign n11994 = ~n11990 & n11993;
  assign n11995 = ~n11057 & n11994;
  assign n11996 = ~n5851 & n11994;
  assign n11997 = ~n11995 & ~n11996;
  assign n11998 =  a[2]  & ~n11997;
  assign n11999 = ~ a[2]  & n11997;
  assign n12000 = ~n11998 & ~n11999;
  assign n12001 = n11989 & n12000;
  assign n12002 = n11469 & n11641;
  assign n12003 = ~n11642 & ~n12002;
  assign n12004 = ~n12001 & n12003;
  assign n12005 = ~n11989 & ~n12000;
  assign n12006 = ~n12004 & ~n12005;
  assign n12007 = ~n1665 & n11727;
  assign n12008 = ~n1877 & n11055;
  assign n12009 = ~n1779 & n11715;
  assign n12010 = ~n12008 & ~n12009;
  assign n12011 = ~n12007 & n12010;
  assign n12012 = ~n11057 & n12011;
  assign n12013 = ~n5328 & n12011;
  assign n12014 = ~n12012 & ~n12013;
  assign n12015 =  a[2]  & ~n12014;
  assign n12016 = ~ a[2]  & n12014;
  assign n12017 = ~n12015 & ~n12016;
  assign n12018 = n12006 & n12017;
  assign n12019 = n11451 & n11643;
  assign n12020 = ~n11644 & ~n12019;
  assign n12021 = ~n12018 & n12020;
  assign n12022 = ~n12006 & ~n12017;
  assign n12023 = ~n12021 & ~n12022;
  assign n12024 = ~n1572 & n11727;
  assign n12025 = ~n1779 & n11055;
  assign n12026 = ~n1665 & n11715;
  assign n12027 = ~n12025 & ~n12026;
  assign n12028 = ~n12024 & n12027;
  assign n12029 = ~n11057 & n12028;
  assign n12030 = ~n5561 & n12028;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 =  a[2]  & ~n12031;
  assign n12033 = ~ a[2]  & n12031;
  assign n12034 = ~n12032 & ~n12033;
  assign n12035 = n12023 & n12034;
  assign n12036 = n11433 & n11645;
  assign n12037 = ~n11646 & ~n12036;
  assign n12038 = ~n12035 & n12037;
  assign n12039 = ~n12023 & ~n12034;
  assign n12040 = ~n12038 & ~n12039;
  assign n12041 = n11647 & ~n11649;
  assign n12042 = ~n11648 & n12041;
  assign n12043 = ~n11651 & ~n12042;
  assign n12044 = ~n12040 & n12043;
  assign n12045 = n12040 & ~n12043;
  assign n12046 = ~n1472 & n11727;
  assign n12047 = ~n1665 & n11055;
  assign n12048 = ~n1572 & n11715;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = ~n12046 & n12049;
  assign n12051 = n5139 & n11057;
  assign n12052 = n12050 & ~n12051;
  assign n12053 = ~ a[2]  & ~n12052;
  assign n12054 =  a[2]  & n12052;
  assign n12055 = ~n12053 & ~n12054;
  assign n12056 = ~n12045 & ~n12055;
  assign n12057 = ~n12044 & ~n12056;
  assign n12058 = n11652 & ~n11654;
  assign n12059 = ~n11653 & n12058;
  assign n12060 = ~n11656 & ~n12059;
  assign n12061 = ~n12057 & n12060;
  assign n12062 = n12057 & ~n12060;
  assign n12063 = ~n1364 & n11727;
  assign n12064 = ~n1572 & n11055;
  assign n12065 = ~n1472 & n11715;
  assign n12066 = ~n12064 & ~n12065;
  assign n12067 = ~n12063 & n12066;
  assign n12068 = n5114 & n11057;
  assign n12069 = n12067 & ~n12068;
  assign n12070 = ~ a[2]  & ~n12069;
  assign n12071 =  a[2]  & n12069;
  assign n12072 = ~n12070 & ~n12071;
  assign n12073 = ~n12062 & ~n12072;
  assign n12074 = ~n12061 & ~n12073;
  assign n12075 = n11787 & ~n12074;
  assign n12076 = ~n11787 & n12074;
  assign n12077 = ~n1235 & n11727;
  assign n12078 = ~n1472 & n11055;
  assign n12079 = ~n1364 & n11715;
  assign n12080 = ~n12078 & ~n12079;
  assign n12081 = ~n12077 & n12080;
  assign n12082 = n4848 & n11057;
  assign n12083 = n12081 & ~n12082;
  assign n12084 = ~ a[2]  & ~n12083;
  assign n12085 =  a[2]  & n12083;
  assign n12086 = ~n12084 & ~n12085;
  assign n12087 = ~n12076 & ~n12086;
  assign n12088 = ~n12075 & ~n12087;
  assign n12089 = ~n1178 & n11727;
  assign n12090 = ~n1364 & n11055;
  assign n12091 = ~n1235 & n11715;
  assign n12092 = ~n12090 & ~n12091;
  assign n12093 = ~n12089 & n12092;
  assign n12094 = ~n11057 & n12093;
  assign n12095 = ~n4861 & n12093;
  assign n12096 = ~n12094 & ~n12095;
  assign n12097 =  a[2]  & ~n12096;
  assign n12098 = ~ a[2]  & n12096;
  assign n12099 = ~n12097 & ~n12098;
  assign n12100 = n12088 & n12099;
  assign n12101 = n11374 & n11661;
  assign n12102 = ~n11662 & ~n12101;
  assign n12103 = ~n12100 & n12102;
  assign n12104 = ~n12088 & ~n12099;
  assign n12105 = ~n12103 & ~n12104;
  assign n12106 = ~n1060 & n11727;
  assign n12107 = ~n1235 & n11055;
  assign n12108 = ~n1178 & n11715;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = ~n12106 & n12109;
  assign n12111 = ~n11057 & n12110;
  assign n12112 = ~n4429 & n12110;
  assign n12113 = ~n12111 & ~n12112;
  assign n12114 =  a[2]  & ~n12113;
  assign n12115 = ~ a[2]  & n12113;
  assign n12116 = ~n12114 & ~n12115;
  assign n12117 = n12105 & n12116;
  assign n12118 = n11356 & n11663;
  assign n12119 = ~n11664 & ~n12118;
  assign n12120 = ~n12117 & n12119;
  assign n12121 = ~n12105 & ~n12116;
  assign n12122 = ~n12120 & ~n12121;
  assign n12123 = ~n958 & n11727;
  assign n12124 = ~n1178 & n11055;
  assign n12125 = ~n1060 & n11715;
  assign n12126 = ~n12124 & ~n12125;
  assign n12127 = ~n12123 & n12126;
  assign n12128 = ~n11057 & n12127;
  assign n12129 = ~n4633 & n12127;
  assign n12130 = ~n12128 & ~n12129;
  assign n12131 =  a[2]  & ~n12130;
  assign n12132 = ~ a[2]  & n12130;
  assign n12133 = ~n12131 & ~n12132;
  assign n12134 = n12122 & n12133;
  assign n12135 = n11338 & n11665;
  assign n12136 = ~n11666 & ~n12135;
  assign n12137 = ~n12134 & n12136;
  assign n12138 = ~n12122 & ~n12133;
  assign n12139 = ~n12137 & ~n12138;
  assign n12140 = n11667 & ~n11669;
  assign n12141 = ~n11668 & n12140;
  assign n12142 = ~n11671 & ~n12141;
  assign n12143 = ~n12139 & n12142;
  assign n12144 = n12139 & ~n12142;
  assign n12145 = ~n867 & n11727;
  assign n12146 = ~n1060 & n11055;
  assign n12147 = ~n958 & n11715;
  assign n12148 = ~n12146 & ~n12147;
  assign n12149 = ~n12145 & n12148;
  assign n12150 = n4204 & n11057;
  assign n12151 = n12149 & ~n12150;
  assign n12152 = ~ a[2]  & ~n12151;
  assign n12153 =  a[2]  & n12151;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = ~n12144 & ~n12154;
  assign n12156 = ~n12143 & ~n12155;
  assign n12157 = n11672 & ~n11674;
  assign n12158 = ~n11673 & n12157;
  assign n12159 = ~n11676 & ~n12158;
  assign n12160 = ~n12156 & n12159;
  assign n12161 = n12156 & ~n12159;
  assign n12162 = ~n710 & n11727;
  assign n12163 = ~n958 & n11055;
  assign n12164 = ~n867 & n11715;
  assign n12165 = ~n12163 & ~n12164;
  assign n12166 = ~n12162 & n12165;
  assign n12167 = n4179 & n11057;
  assign n12168 = n12166 & ~n12167;
  assign n12169 = ~ a[2]  & ~n12168;
  assign n12170 =  a[2]  & n12168;
  assign n12171 = ~n12169 & ~n12170;
  assign n12172 = ~n12161 & ~n12171;
  assign n12173 = ~n12160 & ~n12172;
  assign n12174 = n11785 & ~n12173;
  assign n12175 = ~n11785 & n12173;
  assign n12176 = ~n587 & n11727;
  assign n12177 = ~n867 & n11055;
  assign n12178 = ~n710 & n11715;
  assign n12179 = ~n12177 & ~n12178;
  assign n12180 = ~n12176 & n12179;
  assign n12181 = n3331 & n11057;
  assign n12182 = n12180 & ~n12181;
  assign n12183 = ~ a[2]  & ~n12182;
  assign n12184 =  a[2]  & n12182;
  assign n12185 = ~n12183 & ~n12184;
  assign n12186 = ~n12175 & ~n12185;
  assign n12187 = ~n12174 & ~n12186;
  assign n12188 = ~n392 & n11727;
  assign n12189 = ~n710 & n11055;
  assign n12190 = ~n587 & n11715;
  assign n12191 = ~n12189 & ~n12190;
  assign n12192 = ~n12188 & n12191;
  assign n12193 = ~n11057 & n12192;
  assign n12194 = ~n3347 & n12192;
  assign n12195 = ~n12193 & ~n12194;
  assign n12196 =  a[2]  & ~n12195;
  assign n12197 = ~ a[2]  & n12195;
  assign n12198 = ~n12196 & ~n12197;
  assign n12199 = n12187 & n12198;
  assign n12200 = n11279 & n11681;
  assign n12201 = ~n11682 & ~n12200;
  assign n12202 = ~n12199 & n12201;
  assign n12203 = ~n12187 & ~n12198;
  assign n12204 = ~n12202 & ~n12203;
  assign n12205 = ~n3012 & n11727;
  assign n12206 = ~n587 & n11055;
  assign n12207 = ~n392 & n11715;
  assign n12208 = ~n12206 & ~n12207;
  assign n12209 = ~n12205 & n12208;
  assign n12210 = ~n11057 & n12209;
  assign n12211 = ~n3018 & n12209;
  assign n12212 = ~n12210 & ~n12211;
  assign n12213 =  a[2]  & ~n12212;
  assign n12214 = ~ a[2]  & n12212;
  assign n12215 = ~n12213 & ~n12214;
  assign n12216 = n12204 & n12215;
  assign n12217 = n11261 & n11683;
  assign n12218 = ~n11684 & ~n12217;
  assign n12219 = ~n12216 & n12218;
  assign n12220 = ~n12204 & ~n12215;
  assign n12221 = ~n12219 & ~n12220;
  assign n12222 = ~n3539 & n11727;
  assign n12223 = ~n392 & n11055;
  assign n12224 = ~n3012 & n11715;
  assign n12225 = ~n12223 & ~n12224;
  assign n12226 = ~n12222 & n12225;
  assign n12227 = ~n11057 & n12226;
  assign n12228 = ~n3715 & n12226;
  assign n12229 = ~n12227 & ~n12228;
  assign n12230 =  a[2]  & ~n12229;
  assign n12231 = ~ a[2]  & n12229;
  assign n12232 = ~n12230 & ~n12231;
  assign n12233 = n12221 & n12232;
  assign n12234 = n11243 & n11685;
  assign n12235 = ~n11686 & ~n12234;
  assign n12236 = ~n12233 & n12235;
  assign n12237 = ~n12221 & ~n12232;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = n11687 & ~n11689;
  assign n12240 = ~n11688 & n12239;
  assign n12241 = ~n11691 & ~n12240;
  assign n12242 = ~n12238 & n12241;
  assign n12243 = n12238 & ~n12241;
  assign n12244 = ~n3605 & n11727;
  assign n12245 = ~n3012 & n11055;
  assign n12246 = ~n3539 & n11715;
  assign n12247 = ~n12245 & ~n12246;
  assign n12248 = ~n12244 & n12247;
  assign n12249 = n4084 & n11057;
  assign n12250 = n12248 & ~n12249;
  assign n12251 = ~ a[2]  & ~n12250;
  assign n12252 =  a[2]  & n12250;
  assign n12253 = ~n12251 & ~n12252;
  assign n12254 = ~n12243 & ~n12253;
  assign n12255 = ~n12242 & ~n12254;
  assign n12256 = n11783 & ~n12255;
  assign n12257 = ~n11783 & n12255;
  assign n12258 = ~n3456 & n11727;
  assign n12259 = ~n3539 & n11055;
  assign n12260 = ~n3605 & n11715;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = ~n12258 & n12261;
  assign n12263 = n3627 & n11057;
  assign n12264 = n12262 & ~n12263;
  assign n12265 = ~ a[2]  & ~n12264;
  assign n12266 =  a[2]  & n12264;
  assign n12267 = ~n12265 & ~n12266;
  assign n12268 = ~n12257 & ~n12267;
  assign n12269 = ~n12256 & ~n12268;
  assign n12270 = ~n3805 & n11727;
  assign n12271 = ~n3605 & n11055;
  assign n12272 = ~n3456 & n11715;
  assign n12273 = ~n12271 & ~n12272;
  assign n12274 = ~n12270 & n12273;
  assign n12275 = ~n11057 & n12274;
  assign n12276 = ~n3818 & n12274;
  assign n12277 = ~n12275 & ~n12276;
  assign n12278 =  a[2]  & ~n12277;
  assign n12279 = ~ a[2]  & n12277;
  assign n12280 = ~n12278 & ~n12279;
  assign n12281 = n12269 & n12280;
  assign n12282 = n11198 & n11696;
  assign n12283 = ~n11697 & ~n12282;
  assign n12284 = ~n12281 & n12283;
  assign n12285 = ~n12269 & ~n12280;
  assign n12286 = ~n12284 & ~n12285;
  assign n12287 = n11769 & ~n11781;
  assign n12288 = ~n11780 & ~n11781;
  assign n12289 = ~n12287 & ~n12288;
  assign n12290 = ~n12286 & ~n12289;
  assign n12291 = ~n11781 & ~n12290;
  assign n12292 = ~n11755 & n11766;
  assign n12293 = ~n11767 & ~n12292;
  assign n12294 = ~n12291 & n12293;
  assign n12295 = ~n11767 & ~n12294;
  assign n12296 = ~n11741 & n11752;
  assign n12297 = ~n11753 & ~n12296;
  assign n12298 = ~n12295 & n12297;
  assign n12299 = ~n11753 & ~n12298;
  assign n12300 = ~n11726 & n11738;
  assign n12301 = ~n11739 & ~n12300;
  assign n12302 = ~n12299 & n12301;
  assign n12303 = ~n11739 & ~n12302;
  assign n12304 = ~n11713 & n11723;
  assign n12305 = ~n11724 & ~n12304;
  assign n12306 = ~n12303 & n12305;
  assign n12307 = ~n11724 & ~n12306;
  assign n12308 = n11711 & ~n12307;
  assign n12309 = ~n11709 & ~n12308;
  assign n12310 = n11083 & ~n11086;
  assign n12311 = ~n11087 & ~n12310;
  assign n12312 = ~n12309 & n12311;
  assign n12313 = ~n11087 & ~n12312;
  assign n12314 = n11047 & ~n11049;
  assign n12315 = ~n11050 & ~n12314;
  assign n12316 = ~n12313 & n12315;
  assign n12317 = ~n11050 & ~n12316;
  assign n12318 = n10453 & ~n12317;
  assign n12319 = ~n10451 & ~n12318;
  assign n12320 = n9883 & ~n9886;
  assign n12321 = ~n9887 & ~n12320;
  assign n12322 = ~n12319 & n12321;
  assign n12323 = ~n9887 & ~n12322;
  assign n12324 = n9363 & ~n9365;
  assign n12325 = ~n9366 & ~n12324;
  assign n12326 = ~n12323 & n12325;
  assign n12327 = ~n9366 & ~n12326;
  assign n12328 = n8879 & ~n12327;
  assign n12329 = ~n8877 & ~n12328;
  assign n12330 = n8437 & ~n12329;
  assign n12331 = ~n8435 & ~n12330;
  assign n12332 = n8015 & ~n8017;
  assign n12333 = ~n8018 & ~n12332;
  assign n12334 = ~n12331 & n12333;
  assign n12335 = ~n8018 & ~n12334;
  assign n12336 = n7651 & ~n12335;
  assign n12337 = ~n7649 & ~n12336;
  assign n12338 = n7307 & ~n7310;
  assign n12339 = ~n7311 & ~n12338;
  assign n12340 = ~n12337 & n12339;
  assign n12341 = ~n7311 & ~n12340;
  assign n12342 = n7133 & ~n7135;
  assign n12343 = ~n7136 & ~n12342;
  assign n12344 = ~n12341 & n12343;
  assign n12345 = ~n7136 & ~n12344;
  assign n12346 = n6970 & ~n12345;
  assign n12347 = ~n6968 & ~n12346;
  assign n12348 = n6422 & ~n12347;
  assign n12349 = ~n6420 & ~n12348;
  assign n12350 = n6267 & ~n12349;
  assign n12351 = ~n6265 & ~n12350;
  assign n12352 = n5952 & ~n12351;
  assign n12353 = ~n5950 & ~n12352;
  assign n12354 = n5679 & ~n5681;
  assign n12355 = ~n5682 & ~n12354;
  assign n12356 = ~n12353 & n12355;
  assign n12357 = ~n5682 & ~n12356;
  assign n12358 = n5530 & ~n12357;
  assign n12359 = ~n5528 & ~n12358;
  assign n12360 = n5420 & ~n12359;
  assign n12361 = ~n5418 & ~n12360;
  assign n12362 = n4954 & ~n12361;
  assign n12363 = ~n4952 & ~n12362;
  assign n12364 = n4728 & ~n4730;
  assign n12365 = ~n4731 & ~n12364;
  assign n12366 = ~n12363 & n12365;
  assign n12367 = ~n4731 & ~n12366;
  assign n12368 = n4622 & ~n12367;
  assign n12369 = ~n4622 & n12367;
  assign n12370 = ~n12368 & ~n12369;
  assign n12371 = ~n4621 & ~n12368;
  assign n12372 = ~n4542 & ~n4545;
  assign n12373 = n3457 & ~n3964;
  assign n12374 = ~n3456 & n3542;
  assign n12375 = n3606 & ~n3805;
  assign n12376 = ~n12374 & ~n12375;
  assign n12377 = ~n12373 & n12376;
  assign n12378 = n3368 & n4558;
  assign n12379 = n12377 & ~n12378;
  assign n12380 =  a[29]  & ~n12379;
  assign n12381 =  a[29]  & ~n12380;
  assign n12382 = ~n12379 & ~n12380;
  assign n12383 = ~n12381 & ~n12382;
  assign n12384 = ~n3720 & ~n3724;
  assign n12385 = n288 & n2276;
  assign n12386 = ~n123 & n12385;
  assign n12387 = ~n231 & n12386;
  assign n12388 = ~n495 & n508;
  assign n12389 = ~n367 & n12388;
  assign n12390 = ~n205 & n12389;
  assign n12391 = n2584 & n12390;
  assign n12392 = n12387 & n12391;
  assign n12393 = n2582 & n12392;
  assign n12394 = ~n171 & n12393;
  assign n12395 = ~n121 & n12394;
  assign n12396 = ~n163 & n12395;
  assign n12397 = ~n400 & ~n1203;
  assign n12398 = n1550 & n12397;
  assign n12399 = ~n111 & n12398;
  assign n12400 = ~n289 & n12399;
  assign n12401 = ~n426 & n12400;
  assign n12402 = ~n932 & n12401;
  assign n12403 = ~n470 & n12402;
  assign n12404 = ~n271 & n12403;
  assign n12405 = n533 & n1071;
  assign n12406 = ~n194 & n12405;
  assign n12407 = ~n203 & n12406;
  assign n12408 = ~n147 & n12407;
  assign n12409 = ~n403 & n12408;
  assign n12410 = ~n290 & n2346;
  assign n12411 = ~n452 & n12410;
  assign n12412 = ~n306 & n12411;
  assign n12413 = n1644 & n12412;
  assign n12414 = n12409 & n12413;
  assign n12415 = n1496 & n12414;
  assign n12416 = n2961 & n12415;
  assign n12417 = n811 & n12416;
  assign n12418 = n774 & n12417;
  assign n12419 = n1253 & n12418;
  assign n12420 = n1994 & n12419;
  assign n12421 = n885 & n12420;
  assign n12422 = ~n276 & n12421;
  assign n12423 = ~n847 & n12422;
  assign n12424 = ~n355 & n12423;
  assign n12425 = ~n91 & n12424;
  assign n12426 = ~n424 & n12425;
  assign n12427 = ~n451 & n12426;
  assign n12428 = ~n81 & n12427;
  assign n12429 = ~n142 & ~n301;
  assign n12430 = ~n564 & n12429;
  assign n12431 = ~n633 & n12430;
  assign n12432 = n253 & n722;
  assign n12433 = n1158 & n12432;
  assign n12434 = n12431 & n12433;
  assign n12435 = n12428 & n12434;
  assign n12436 = n12404 & n12435;
  assign n12437 = n6769 & n12436;
  assign n12438 = n12396 & n12437;
  assign n12439 = n3163 & n12438;
  assign n12440 = ~n1306 & n12439;
  assign n12441 = ~n232 & n12440;
  assign n12442 = ~n571 & n12441;
  assign n12443 = ~n656 & n12442;
  assign n12444 = ~n357 & n12443;
  assign n12445 = ~n371 & n12444;
  assign n12446 = ~n119 & n12445;
  assign n12447 = ~n569 & n12446;
  assign n12448 = ~n429 & n12447;
  assign n12449 = ~n3702 & ~n12448;
  assign n12450 = n3702 & n12448;
  assign n12451 = ~n12449 & ~n12450;
  assign n12452 = ~ a[23]  & n12451;
  assign n12453 = ~ a[23]  & ~n12452;
  assign n12454 = ~n12449 & ~n12452;
  assign n12455 = ~n12450 & n12454;
  assign n12456 = ~n12453 & ~n12455;
  assign n12457 = n3020 & ~n3605;
  assign n12458 = n3028 & ~n3539;
  assign n12459 = ~n3012 & n3023;
  assign n12460 = n75 & n4084;
  assign n12461 = ~n12459 & ~n12460;
  assign n12462 = ~n12458 & n12461;
  assign n12463 = ~n12457 & n12462;
  assign n12464 = ~n12456 & ~n12463;
  assign n12465 = n12456 & n12463;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = ~n3708 & n12466;
  assign n12468 = n3708 & ~n12466;
  assign n12469 = ~n12467 & ~n12468;
  assign n12470 = ~n12384 & n12469;
  assign n12471 = n12384 & ~n12469;
  assign n12472 = ~n12470 & ~n12471;
  assign n12473 = ~n12383 & n12472;
  assign n12474 = n12472 & ~n12473;
  assign n12475 = ~n12383 & ~n12473;
  assign n12476 = ~n12474 & ~n12475;
  assign n12477 = ~n3825 & ~n4074;
  assign n12478 = n3884 & ~n4515;
  assign n12479 = n3967 & ~n4045;
  assign n12480 = ~n3877 & n4046;
  assign n12481 = ~n12479 & ~n12480;
  assign n12482 = ~n12478 & n12481;
  assign n12483 = ~n4050 & n12482;
  assign n12484 = ~n4715 & n12482;
  assign n12485 = ~n12483 & ~n12484;
  assign n12486 =  a[26]  & ~n12485;
  assign n12487 = ~ a[26]  & n12485;
  assign n12488 = ~n12486 & ~n12487;
  assign n12489 = ~n12477 & ~n12488;
  assign n12490 = ~n12477 & ~n12489;
  assign n12491 = ~n12488 & ~n12489;
  assign n12492 = ~n12490 & ~n12491;
  assign n12493 = ~n12476 & ~n12492;
  assign n12494 = n12476 & ~n12491;
  assign n12495 = ~n12490 & n12494;
  assign n12496 = ~n12493 & ~n12495;
  assign n12497 = ~n12372 & n12496;
  assign n12498 = n12372 & ~n12496;
  assign n12499 = ~n12497 & ~n12498;
  assign n12500 = ~n12371 & n12499;
  assign n12501 = n12371 & ~n12499;
  assign n12502 = ~n12500 & ~n12501;
  assign n12503 = n12370 & n12502;
  assign n12504 = n12363 & ~n12365;
  assign n12505 = ~n12366 & ~n12504;
  assign n12506 = n12370 & n12505;
  assign n12507 = ~n4954 & n12361;
  assign n12508 = ~n12362 & ~n12507;
  assign n12509 = n12505 & n12508;
  assign n12510 = ~n5530 & n12357;
  assign n12511 = ~n12358 & ~n12510;
  assign n12512 = ~n5420 & n12359;
  assign n12513 = ~n12360 & ~n12512;
  assign n12514 = n12511 & n12513;
  assign n12515 = n12353 & ~n12355;
  assign n12516 = ~n12356 & ~n12515;
  assign n12517 = n12511 & n12516;
  assign n12518 = ~n5952 & n12351;
  assign n12519 = ~n12352 & ~n12518;
  assign n12520 = n12516 & n12519;
  assign n12521 = ~n6267 & n12349;
  assign n12522 = ~n12350 & ~n12521;
  assign n12523 = n12519 & n12522;
  assign n12524 = ~n6422 & n12347;
  assign n12525 = ~n12348 & ~n12524;
  assign n12526 = n12522 & n12525;
  assign n12527 = ~n6970 & n12345;
  assign n12528 = ~n12346 & ~n12527;
  assign n12529 = n12525 & n12528;
  assign n12530 = n12341 & ~n12343;
  assign n12531 = ~n12344 & ~n12530;
  assign n12532 = n12528 & n12531;
  assign n12533 = n12337 & ~n12339;
  assign n12534 = ~n12340 & ~n12533;
  assign n12535 = n12531 & n12534;
  assign n12536 = ~n7651 & n12335;
  assign n12537 = ~n12336 & ~n12536;
  assign n12538 = n12534 & n12537;
  assign n12539 = n12331 & ~n12333;
  assign n12540 = ~n12334 & ~n12539;
  assign n12541 = n12537 & n12540;
  assign n12542 = ~n8437 & n12329;
  assign n12543 = ~n12330 & ~n12542;
  assign n12544 = n12540 & n12543;
  assign n12545 = ~n8879 & n12327;
  assign n12546 = ~n12328 & ~n12545;
  assign n12547 = n12543 & n12546;
  assign n12548 = n12323 & ~n12325;
  assign n12549 = ~n12326 & ~n12548;
  assign n12550 = n12546 & n12549;
  assign n12551 = n12319 & ~n12321;
  assign n12552 = ~n12322 & ~n12551;
  assign n12553 = n12549 & n12552;
  assign n12554 = ~n10453 & n12317;
  assign n12555 = ~n12318 & ~n12554;
  assign n12556 = n12552 & n12555;
  assign n12557 = n12313 & ~n12315;
  assign n12558 = ~n12316 & ~n12557;
  assign n12559 = n12555 & n12558;
  assign n12560 = n12309 & ~n12311;
  assign n12561 = ~n12312 & ~n12560;
  assign n12562 = n12558 & n12561;
  assign n12563 = ~n11711 & n12307;
  assign n12564 = ~n12308 & ~n12563;
  assign n12565 = n12561 & n12564;
  assign n12566 = n12303 & ~n12305;
  assign n12567 = ~n12306 & ~n12566;
  assign n12568 = n12564 & n12567;
  assign n12569 = ~n12564 & ~n12567;
  assign n12570 = n12299 & ~n12301;
  assign n12571 = ~n12302 & ~n12570;
  assign n12572 = n12567 & n12571;
  assign n12573 = n12295 & ~n12297;
  assign n12574 = ~n12298 & ~n12573;
  assign n12575 = n12571 & n12574;
  assign n12576 = n12291 & ~n12293;
  assign n12577 = ~n12294 & ~n12576;
  assign n12578 = n12574 & n12577;
  assign n12579 = ~n12286 & ~n12290;
  assign n12580 = ~n12289 & ~n12290;
  assign n12581 = ~n12579 & ~n12580;
  assign n12582 = n12577 & ~n12581;
  assign n12583 = ~n12574 & n12582;
  assign n12584 = ~n12578 & ~n12583;
  assign n12585 = ~n12571 & ~n12574;
  assign n12586 = ~n12575 & ~n12585;
  assign n12587 = ~n12584 & n12586;
  assign n12588 = ~n12575 & ~n12587;
  assign n12589 = ~n12567 & ~n12571;
  assign n12590 = ~n12572 & ~n12589;
  assign n12591 = ~n12588 & n12590;
  assign n12592 = ~n12572 & ~n12591;
  assign n12593 = ~n12568 & ~n12592;
  assign n12594 = ~n12569 & n12593;
  assign n12595 = ~n12568 & ~n12594;
  assign n12596 = ~n12561 & ~n12564;
  assign n12597 = ~n12595 & ~n12596;
  assign n12598 = ~n12565 & n12597;
  assign n12599 = ~n12565 & ~n12598;
  assign n12600 = ~n12558 & ~n12561;
  assign n12601 = ~n12562 & ~n12600;
  assign n12602 = ~n12599 & n12601;
  assign n12603 = ~n12562 & ~n12602;
  assign n12604 = ~n12555 & ~n12558;
  assign n12605 = ~n12603 & ~n12604;
  assign n12606 = ~n12559 & n12605;
  assign n12607 = ~n12559 & ~n12606;
  assign n12608 = ~n12552 & ~n12555;
  assign n12609 = ~n12607 & ~n12608;
  assign n12610 = ~n12556 & n12609;
  assign n12611 = ~n12556 & ~n12610;
  assign n12612 = ~n12549 & ~n12552;
  assign n12613 = ~n12553 & ~n12612;
  assign n12614 = ~n12611 & n12613;
  assign n12615 = ~n12553 & ~n12614;
  assign n12616 = ~n12546 & ~n12549;
  assign n12617 = ~n12615 & ~n12616;
  assign n12618 = ~n12550 & n12617;
  assign n12619 = ~n12550 & ~n12618;
  assign n12620 = ~n12543 & ~n12546;
  assign n12621 = ~n12547 & ~n12620;
  assign n12622 = ~n12619 & n12621;
  assign n12623 = ~n12547 & ~n12622;
  assign n12624 = ~n12540 & ~n12543;
  assign n12625 = ~n12623 & ~n12624;
  assign n12626 = ~n12544 & n12625;
  assign n12627 = ~n12544 & ~n12626;
  assign n12628 = ~n12537 & ~n12540;
  assign n12629 = ~n12627 & ~n12628;
  assign n12630 = ~n12541 & n12629;
  assign n12631 = ~n12541 & ~n12630;
  assign n12632 = ~n12534 & ~n12537;
  assign n12633 = ~n12631 & ~n12632;
  assign n12634 = ~n12538 & n12633;
  assign n12635 = ~n12538 & ~n12634;
  assign n12636 = ~n12531 & ~n12534;
  assign n12637 = ~n12535 & ~n12636;
  assign n12638 = ~n12635 & n12637;
  assign n12639 = ~n12535 & ~n12638;
  assign n12640 = ~n12528 & ~n12531;
  assign n12641 = ~n12639 & ~n12640;
  assign n12642 = ~n12532 & n12641;
  assign n12643 = ~n12532 & ~n12642;
  assign n12644 = ~n12525 & ~n12528;
  assign n12645 = ~n12529 & ~n12644;
  assign n12646 = ~n12643 & n12645;
  assign n12647 = ~n12529 & ~n12646;
  assign n12648 = ~n12522 & ~n12525;
  assign n12649 = ~n12526 & ~n12648;
  assign n12650 = ~n12647 & n12649;
  assign n12651 = ~n12526 & ~n12650;
  assign n12652 = ~n12519 & ~n12522;
  assign n12653 = ~n12523 & ~n12652;
  assign n12654 = ~n12651 & n12653;
  assign n12655 = ~n12523 & ~n12654;
  assign n12656 = ~n12516 & ~n12519;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = ~n12520 & n12657;
  assign n12659 = ~n12520 & ~n12658;
  assign n12660 = ~n12511 & ~n12516;
  assign n12661 = ~n12659 & ~n12660;
  assign n12662 = ~n12517 & n12661;
  assign n12663 = ~n12517 & ~n12662;
  assign n12664 = ~n12511 & ~n12513;
  assign n12665 = ~n12514 & ~n12664;
  assign n12666 = ~n12663 & n12665;
  assign n12667 = ~n12514 & ~n12666;
  assign n12668 = ~n12508 & ~n12513;
  assign n12669 = n12508 & n12513;
  assign n12670 = ~n12668 & ~n12669;
  assign n12671 = ~n12667 & n12670;
  assign n12672 = ~n12669 & ~n12671;
  assign n12673 = ~n12505 & ~n12508;
  assign n12674 = ~n12672 & ~n12673;
  assign n12675 = ~n12509 & n12674;
  assign n12676 = ~n12509 & ~n12675;
  assign n12677 = ~n12370 & ~n12505;
  assign n12678 = ~n12676 & ~n12677;
  assign n12679 = ~n12506 & n12678;
  assign n12680 = ~n12506 & ~n12679;
  assign n12681 = ~n12370 & ~n12502;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = ~n12503 & n12682;
  assign n12684 = ~n12503 & ~n12683;
  assign n12685 = ~n12497 & ~n12500;
  assign n12686 = ~n12489 & ~n12493;
  assign n12687 = ~n3877 & n3967;
  assign n12688 = n4046 & ~n4515;
  assign n12689 = ~n12687 & ~n12688;
  assign n12690 = n4050 & n4609;
  assign n12691 = n12689 & ~n12690;
  assign n12692 =  a[26]  & ~n12691;
  assign n12693 = ~n12691 & ~n12692;
  assign n12694 =  a[26]  & ~n12692;
  assign n12695 = ~n12693 & ~n12694;
  assign n12696 = ~n12470 & ~n12473;
  assign n12697 = n75 & n3627;
  assign n12698 = n3020 & ~n3456;
  assign n12699 = n3023 & ~n3539;
  assign n12700 = n3028 & ~n3605;
  assign n12701 = ~n12699 & ~n12700;
  assign n12702 = ~n12698 & n12701;
  assign n12703 = ~n12697 & n12702;
  assign n12704 = ~n169 & ~n194;
  assign n12705 = ~n803 & n12704;
  assign n12706 = ~n1101 & n12705;
  assign n12707 = ~n419 & n12706;
  assign n12708 = ~n394 & n12707;
  assign n12709 = ~n657 & n12708;
  assign n12710 = ~n161 & n12709;
  assign n12711 = ~n232 & ~n393;
  assign n12712 = ~n201 & n12711;
  assign n12713 = n2361 & n12712;
  assign n12714 = n1879 & n12713;
  assign n12715 = n6054 & n12714;
  assign n12716 = n5806 & n12715;
  assign n12717 = n1549 & n12716;
  assign n12718 = n2507 & n12717;
  assign n12719 = n1577 & n12718;
  assign n12720 = n2573 & n12719;
  assign n12721 = n12710 & n12720;
  assign n12722 = n120 & n12721;
  assign n12723 = n4786 & n12722;
  assign n12724 = n356 & n12723;
  assign n12725 = n116 & n12724;
  assign n12726 = ~n154 & n12725;
  assign n12727 = ~n715 & n12726;
  assign n12728 = ~n102 & n12727;
  assign n12729 = ~n277 & n12728;
  assign n12730 = ~n270 & n12729;
  assign n12731 = ~n12454 & n12730;
  assign n12732 = n12454 & ~n12730;
  assign n12733 = ~n12731 & ~n12732;
  assign n12734 = ~n12703 & n12733;
  assign n12735 = ~n12703 & ~n12734;
  assign n12736 = n12733 & ~n12734;
  assign n12737 = ~n12735 & ~n12736;
  assign n12738 = ~n12464 & ~n12467;
  assign n12739 = n12737 & n12738;
  assign n12740 = ~n12737 & ~n12738;
  assign n12741 = ~n12739 & ~n12740;
  assign n12742 = n3457 & ~n4045;
  assign n12743 = n3542 & ~n3805;
  assign n12744 = n3606 & ~n3964;
  assign n12745 = ~n12743 & ~n12744;
  assign n12746 = ~n12742 & n12745;
  assign n12747 = ~n3368 & n12746;
  assign n12748 = ~n4477 & n12746;
  assign n12749 = ~n12747 & ~n12748;
  assign n12750 =  a[29]  & ~n12749;
  assign n12751 = ~ a[29]  & n12749;
  assign n12752 = ~n12750 & ~n12751;
  assign n12753 = n12741 & ~n12752;
  assign n12754 = ~n12741 & n12752;
  assign n12755 = ~n12753 & ~n12754;
  assign n12756 = ~n12696 & n12755;
  assign n12757 = ~n12696 & ~n12756;
  assign n12758 = n12755 & ~n12756;
  assign n12759 = ~n12757 & ~n12758;
  assign n12760 = ~n12695 & ~n12759;
  assign n12761 = n12695 & ~n12758;
  assign n12762 = ~n12757 & n12761;
  assign n12763 = ~n12760 & ~n12762;
  assign n12764 = ~n12686 & n12763;
  assign n12765 = n12686 & ~n12763;
  assign n12766 = ~n12764 & ~n12765;
  assign n12767 = ~n12685 & n12766;
  assign n12768 = n12685 & ~n12766;
  assign n12769 = ~n12767 & ~n12768;
  assign n12770 = ~n12502 & ~n12769;
  assign n12771 = n12502 & n12769;
  assign n12772 = ~n12770 & ~n12771;
  assign n12773 = ~n12684 & n12772;
  assign n12774 = ~n12771 & ~n12773;
  assign n12775 = ~n12764 & ~n12767;
  assign n12776 = ~n12756 & ~n12760;
  assign n12777 = n75 & n3818;
  assign n12778 = n3020 & ~n3805;
  assign n12779 = n3023 & ~n3605;
  assign n12780 = n3028 & ~n3456;
  assign n12781 = ~n12779 & ~n12780;
  assign n12782 = ~n12778 & n12781;
  assign n12783 = ~n12777 & n12782;
  assign n12784 = ~n224 & ~n305;
  assign n12785 = ~n714 & n12784;
  assign n12786 = n653 & n12785;
  assign n12787 = n2573 & n12786;
  assign n12788 = n2582 & n12787;
  assign n12789 = ~n276 & n12788;
  assign n12790 = ~n460 & n12789;
  assign n12791 = ~n932 & n12790;
  assign n12792 = ~n273 & n12791;
  assign n12793 = ~n225 & n12792;
  assign n12794 = ~n712 & n12793;
  assign n12795 = ~n231 & n12794;
  assign n12796 = n561 & n5808;
  assign n12797 = n1476 & n12796;
  assign n12798 = n968 & n12797;
  assign n12799 = n2170 & n12798;
  assign n12800 = n282 & n12799;
  assign n12801 = n1247 & n12800;
  assign n12802 = ~n206 & n12801;
  assign n12803 = ~n673 & n12802;
  assign n12804 = ~n531 & n12803;
  assign n12805 = ~n1104 & n12804;
  assign n12806 = ~n462 & ~n667;
  assign n12807 = ~n151 & n12806;
  assign n12808 = ~n1062 & n12807;
  assign n12809 = ~n451 & n12808;
  assign n12810 = ~n125 & n12809;
  assign n12811 = ~n403 & ~n506;
  assign n12812 = ~n601 & n12811;
  assign n12813 = n1527 & n12812;
  assign n12814 = n12810 & n12813;
  assign n12815 = n12805 & n12814;
  assign n12816 = n4794 & n12815;
  assign n12817 = n202 & n12816;
  assign n12818 = ~n190 & n12817;
  assign n12819 = ~n255 & n12818;
  assign n12820 = ~n239 & n12819;
  assign n12821 = ~n121 & n12820;
  assign n12822 = ~n402 & n12821;
  assign n12823 = ~n287 & n12822;
  assign n12824 = ~n302 & n12823;
  assign n12825 = ~n243 & n12824;
  assign n12826 = ~n519 & n12825;
  assign n12827 = ~n271 & n12826;
  assign n12828 = ~n429 & n12827;
  assign n12829 = ~n334 & ~n435;
  assign n12830 = ~n252 & n12829;
  assign n12831 = n3827 & n12830;
  assign n12832 = n6084 & n12831;
  assign n12833 = n12828 & n12832;
  assign n12834 = n12795 & n12833;
  assign n12835 = n1479 & n12834;
  assign n12836 = n159 & n12835;
  assign n12837 = n1667 & n12836;
  assign n12838 = n570 & n12837;
  assign n12839 = ~n284 & n12838;
  assign n12840 = ~n191 & n12839;
  assign n12841 = ~n452 & n12840;
  assign n12842 = ~n474 & n12841;
  assign n12843 = ~n12730 & n12842;
  assign n12844 = n12730 & ~n12842;
  assign n12845 = ~n12783 & ~n12844;
  assign n12846 = ~n12843 & n12845;
  assign n12847 = ~n12783 & ~n12846;
  assign n12848 = ~n12844 & ~n12846;
  assign n12849 = ~n12843 & n12848;
  assign n12850 = ~n12847 & ~n12849;
  assign n12851 = ~n12731 & ~n12734;
  assign n12852 = n12850 & n12851;
  assign n12853 = ~n12850 & ~n12851;
  assign n12854 = ~n12852 & ~n12853;
  assign n12855 = ~n12740 & ~n12753;
  assign n12856 = n12854 & ~n12855;
  assign n12857 = ~n12854 & n12855;
  assign n12858 = ~n12856 & ~n12857;
  assign n12859 = n4050 & n4522;
  assign n12860 = n3967 & ~n4515;
  assign n12861 = ~n12859 & ~n12860;
  assign n12862 =  a[26]  & ~n12861;
  assign n12863 = ~n12861 & ~n12862;
  assign n12864 =  a[26]  & ~n12862;
  assign n12865 = ~n12863 & ~n12864;
  assign n12866 = n3457 & ~n3877;
  assign n12867 = n3542 & ~n3964;
  assign n12868 = n3606 & ~n4045;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = ~n12866 & n12869;
  assign n12871 = n3368 & n4067;
  assign n12872 = n12870 & ~n12871;
  assign n12873 =  a[29]  & ~n12872;
  assign n12874 =  a[29]  & ~n12873;
  assign n12875 = ~n12872 & ~n12873;
  assign n12876 = ~n12874 & ~n12875;
  assign n12877 = ~n12865 & ~n12876;
  assign n12878 = ~n12865 & ~n12877;
  assign n12879 = ~n12876 & ~n12877;
  assign n12880 = ~n12878 & ~n12879;
  assign n12881 = n12858 & ~n12880;
  assign n12882 = ~n12858 & n12880;
  assign n12883 = ~n12881 & ~n12882;
  assign n12884 = ~n12776 & n12883;
  assign n12885 = n12776 & ~n12883;
  assign n12886 = ~n12884 & ~n12885;
  assign n12887 = ~n12775 & n12886;
  assign n12888 = n12775 & ~n12886;
  assign n12889 = ~n12887 & ~n12888;
  assign n12890 = ~n12769 & ~n12889;
  assign n12891 = n12769 & n12889;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = ~n12774 & n12892;
  assign n12894 = n12774 & ~n12892;
  assign n12895 = ~n12893 & ~n12894;
  assign n12896 = n75 & n12895;
  assign n12897 = n3020 & n12889;
  assign n12898 = n3023 & n12502;
  assign n12899 = n3028 & n12769;
  assign n12900 = ~n12898 & ~n12899;
  assign n12901 = ~n12897 & n12900;
  assign n12902 = ~n12896 & n12901;
  assign n12903 = ~n276 & ~n667;
  assign n12904 = ~n190 & n12903;
  assign n12905 = ~n1101 & n12904;
  assign n12906 = ~n396 & n12905;
  assign n12907 = ~n453 & n12906;
  assign n12908 = ~n422 & n12907;
  assign n12909 = ~n132 & n12908;
  assign n12910 = n230 & ~n306;
  assign n12911 = ~n272 & n12910;
  assign n12912 = n1611 & n4327;
  assign n12913 = n12911 & n12912;
  assign n12914 = ~n155 & n12913;
  assign n12915 = ~n402 & n12914;
  assign n12916 = ~n1104 & n12915;
  assign n12917 = ~n883 & n12916;
  assign n12918 = ~n337 & n12917;
  assign n12919 = ~n188 & n12918;
  assign n12920 = ~n239 & n2092;
  assign n12921 = ~n825 & n12920;
  assign n12922 = ~n601 & n12921;
  assign n12923 = ~n567 & n12922;
  assign n12924 = ~n293 & n12923;
  assign n12925 = n1994 & n6520;
  assign n12926 = n1782 & n12925;
  assign n12927 = ~n111 & n12926;
  assign n12928 = ~n242 & n12927;
  assign n12929 = ~n327 & n12928;
  assign n12930 = ~n147 & n12929;
  assign n12931 = ~n395 & n12930;
  assign n12932 = ~n86 & n12931;
  assign n12933 = n640 & n5040;
  assign n12934 = n12932 & n12933;
  assign n12935 = n12924 & n12934;
  assign n12936 = n2443 & n12935;
  assign n12937 = ~n136 & n12936;
  assign n12938 = ~n886 & n12937;
  assign n12939 = ~n358 & n12938;
  assign n12940 = ~n355 & ~n1011;
  assign n12941 = ~n171 & n12940;
  assign n12942 = n373 & n12941;
  assign n12943 = n1237 & n12942;
  assign n12944 = ~n564 & n12943;
  assign n12945 = n638 & n2230;
  assign n12946 = n1249 & n12945;
  assign n12947 = n2468 & n12946;
  assign n12948 = n12944 & n12947;
  assign n12949 = n12939 & n12948;
  assign n12950 = n2623 & n12949;
  assign n12951 = n12919 & n12950;
  assign n12952 = n12909 & n12951;
  assign n12953 = n1129 & n12952;
  assign n12954 = n4295 & n12953;
  assign n12955 = ~n330 & n12954;
  assign n12956 = ~n254 & n12955;
  assign n12957 = ~n292 & n12956;
  assign n12958 = ~n91 & n12957;
  assign n12959 = n2684 & n3438;
  assign n12960 = n530 & n12959;
  assign n12961 = n1925 & n12960;
  assign n12962 = n789 & n12961;
  assign n12963 = n1254 & n12962;
  assign n12964 = n1827 & n12963;
  assign n12965 = n1161 & n12964;
  assign n12966 = ~n847 & n12965;
  assign n12967 = ~n619 & n12966;
  assign n12968 = ~n155 & n12967;
  assign n12969 = ~n637 & n12968;
  assign n12970 = ~n980 & n12969;
  assign n12971 = ~n394 & n12970;
  assign n12972 = ~n225 & n12971;
  assign n12973 = ~n332 & n12972;
  assign n12974 = ~n281 & ~n426;
  assign n12975 = ~n189 & n12974;
  assign n12976 = ~n461 & n12975;
  assign n12977 = ~n231 & n12976;
  assign n12978 = n3985 & n4334;
  assign n12979 = n12977 & n12978;
  assign n12980 = n1216 & n12979;
  assign n12981 = n5224 & n12980;
  assign n12982 = n1969 & n12981;
  assign n12983 = n12973 & n12982;
  assign n12984 = n1523 & n12983;
  assign n12985 = n2633 & n12984;
  assign n12986 = n1825 & n12985;
  assign n12987 = n1252 & n12986;
  assign n12988 = ~n242 & n12987;
  assign n12989 = ~n355 & n12988;
  assign n12990 = ~n495 & n12989;
  assign n12991 = ~n246 & n12990;
  assign n12992 = n6706 & n12991;
  assign n12993 = ~n375 & n12992;
  assign n12994 = ~n237 & n12993;
  assign n12995 = ~n564 & n12994;
  assign n12996 = n12958 & ~n12995;
  assign n12997 = ~n12958 & n12995;
  assign n12998 = n12684 & ~n12772;
  assign n12999 = ~n12773 & ~n12998;
  assign n13000 = n75 & n12999;
  assign n13001 = n3020 & n12769;
  assign n13002 = n3023 & n12370;
  assign n13003 = n3028 & n12502;
  assign n13004 = ~n13002 & ~n13003;
  assign n13005 = ~n13001 & n13004;
  assign n13006 = ~n13000 & n13005;
  assign n13007 = ~n12996 & ~n13006;
  assign n13008 = ~n12997 & n13007;
  assign n13009 = ~n12996 & ~n13008;
  assign n13010 = ~n169 & n238;
  assign n13011 = ~n514 & n13010;
  assign n13012 = ~n119 & n13011;
  assign n13013 = ~n353 & ~n847;
  assign n13014 = ~n326 & n13013;
  assign n13015 = ~n419 & ~n689;
  assign n13016 = ~n493 & n13015;
  assign n13017 = n13014 & n13016;
  assign n13018 = n1693 & n13017;
  assign n13019 = n13012 & n13018;
  assign n13020 = n12795 & n13019;
  assign n13021 = n1511 & n13020;
  assign n13022 = n2782 & n13021;
  assign n13023 = n2507 & n13022;
  assign n13024 = n1827 & n13023;
  assign n13025 = n1248 & n13024;
  assign n13026 = ~n301 & n13025;
  assign n13027 = ~n278 & n13026;
  assign n13028 = ~n115 & n13027;
  assign n13029 = ~n91 & n13028;
  assign n13030 = ~n504 & n13029;
  assign n13031 = ~n436 & n13030;
  assign n13032 = n1556 & n4151;
  assign n13033 = n897 & n13032;
  assign n13034 = n591 & n13033;
  assign n13035 = ~n656 & n13034;
  assign n13036 = ~n594 & n13035;
  assign n13037 = ~n417 & n13036;
  assign n13038 = ~n527 & n13037;
  assign n13039 = ~n165 & n13038;
  assign n13040 = ~n672 & n13039;
  assign n13041 = ~n293 & n13040;
  assign n13042 = n2020 & n6664;
  assign n13043 = n593 & n13042;
  assign n13044 = n6607 & n13043;
  assign n13045 = n12828 & n13044;
  assign n13046 = n13041 & n13045;
  assign n13047 = n1521 & n13046;
  assign n13048 = n13031 & n13047;
  assign n13049 = n1029 & n13048;
  assign n13050 = n291 & n13049;
  assign n13051 = n1139 & n13050;
  assign n13052 = n826 & n13051;
  assign n13053 = n1389 & n13052;
  assign n13054 = n341 & n13053;
  assign n13055 = ~n1102 & n13054;
  assign n13056 = ~n1127 & n13055;
  assign n13057 = n3831 & n13056;
  assign n13058 = n193 & n13057;
  assign n13059 = ~n452 & n13058;
  assign n13060 = n1255 & n1781;
  assign n13061 = n3984 & n13060;
  assign n13062 = ~n589 & n13061;
  assign n13063 = ~n449 & n13062;
  assign n13064 = n2265 & n3906;
  assign n13065 = n3580 & n13064;
  assign n13066 = n5233 & n13065;
  assign n13067 = n4017 & n13066;
  assign n13068 = n13063 & n13067;
  assign n13069 = n4502 & n13068;
  assign n13070 = n3848 & n13069;
  assign n13071 = n2738 & n13070;
  assign n13072 = n2583 & n13071;
  assign n13073 = ~n242 & n13072;
  assign n13074 = ~n518 & n13073;
  assign n13075 = n3569 & n3906;
  assign n13076 = n3832 & n4034;
  assign n13077 = n13075 & n13076;
  assign n13078 = n3869 & n13077;
  assign n13079 = ~n328 & n13078;
  assign n13080 = ~n536 & n13079;
  assign n13081 = ~n567 & n13080;
  assign n13082 = n13074 & n13081;
  assign n13083 = ~n13059 & n13082;
  assign n13084 = n3570 & n3832;
  assign n13085 = n539 & n13084;
  assign n13086 = n968 & n13085;
  assign n13087 = ~n453 & n13086;
  assign n13088 = n3949 & n13087;
  assign n13089 = n3856 & n13088;
  assign n13090 = n4493 & n13089;
  assign n13091 = n665 & n13090;
  assign n13092 = n1761 & n13091;
  assign n13093 = ~n601 & n13092;
  assign n13094 = ~n673 & n13093;
  assign n13095 = ~n99 & n13094;
  assign n13096 = n13074 & ~n13095;
  assign n13097 = ~n13074 & n13095;
  assign n13098 = n75 & n4522;
  assign n13099 = n3023 & ~n4515;
  assign n13100 = ~n13098 & ~n13099;
  assign n13101 = ~n13096 & ~n13100;
  assign n13102 = ~n13097 & n13101;
  assign n13103 = ~n13096 & ~n13102;
  assign n13104 = ~n13074 & ~n13081;
  assign n13105 = ~n13082 & ~n13104;
  assign n13106 = ~n13103 & ~n13105;
  assign n13107 = ~n13103 & ~n13106;
  assign n13108 = ~n13105 & ~n13106;
  assign n13109 = ~n13107 & ~n13108;
  assign n13110 = ~n13100 & ~n13102;
  assign n13111 = ~n13097 & n13103;
  assign n13112 = ~n13110 & ~n13111;
  assign n13113 = ~n283 & ~n1306;
  assign n13114 = ~n249 & n13113;
  assign n13115 = n12397 & n13114;
  assign n13116 = n4216 & n13115;
  assign n13117 = n1916 & n13116;
  assign n13118 = ~n305 & n13117;
  assign n13119 = ~n403 & n13118;
  assign n13120 = ~n246 & n13119;
  assign n13121 = ~n519 & n13120;
  assign n13122 = ~n125 & n13121;
  assign n13123 = ~n293 & n13122;
  assign n13124 = n530 & n3570;
  assign n13125 = n2740 & n13124;
  assign n13126 = ~n232 & n13125;
  assign n13127 = ~n289 & n13126;
  assign n13128 = ~n149 & n13127;
  assign n13129 = ~n226 & n13128;
  assign n13130 = ~n490 & n13129;
  assign n13131 = ~n496 & n13130;
  assign n13132 = ~n157 & n13131;
  assign n13133 = ~n623 & n13132;
  assign n13134 = ~n86 & n13133;
  assign n13135 = ~n771 & n13134;
  assign n13136 = ~n167 & n13135;
  assign n13137 = ~n165 & n13136;
  assign n13138 = ~n158 & n13137;
  assign n13139 = n1163 & n2544;
  assign n13140 = n13138 & n13139;
  assign n13141 = n1735 & n13140;
  assign n13142 = n1202 & n13141;
  assign n13143 = n13123 & n13142;
  assign n13144 = n5085 & n13143;
  assign n13145 = n2635 & n13144;
  assign n13146 = n1366 & n13145;
  assign n13147 = n730 & n13146;
  assign n13148 = n1252 & n13147;
  assign n13149 = n2466 & n13148;
  assign n13150 = n978 & n13149;
  assign n13151 = ~n123 & n13150;
  assign n13152 = ~n847 & n13151;
  assign n13153 = ~n284 & n13152;
  assign n13154 = ~n367 & n13153;
  assign n13155 = ~n292 & n13154;
  assign n13156 = ~n274 & n13155;
  assign n13157 = ~n525 & n13156;
  assign n13158 = ~n672 & n13157;
  assign n13159 = n3929 & n5064;
  assign n13160 = n885 & n13159;
  assign n13161 = ~n144 & n13160;
  assign n13162 = n1425 & n1740;
  assign n13163 = n1249 & n13162;
  assign n13164 = n13161 & n13163;
  assign n13165 = n13087 & n13164;
  assign n13166 = n3947 & n13165;
  assign n13167 = n13063 & n13166;
  assign n13168 = n4009 & n13167;
  assign n13169 = n1046 & n13168;
  assign n13170 = ~n567 & n13169;
  assign n13171 = ~n525 & n13170;
  assign n13172 = ~n293 & n13171;
  assign n13173 = ~n13158 & ~n13172;
  assign n13174 = n13158 & n13172;
  assign n13175 = ~n13173 & ~n13174;
  assign n13176 = ~ a[29]  & n13175;
  assign n13177 = ~n13173 & ~n13176;
  assign n13178 = n13074 & ~n13177;
  assign n13179 = n75 & n4609;
  assign n13180 = n3023 & ~n3877;
  assign n13181 = n3028 & ~n4515;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = ~n13179 & n13182;
  assign n13184 = ~n13074 & n13177;
  assign n13185 = ~n13178 & ~n13184;
  assign n13186 = ~n13183 & n13185;
  assign n13187 = ~n13178 & ~n13186;
  assign n13188 = ~n13112 & ~n13187;
  assign n13189 = n13112 & n13187;
  assign n13190 = ~n13188 & ~n13189;
  assign n13191 = ~n13183 & ~n13186;
  assign n13192 = n13185 & ~n13186;
  assign n13193 = ~n13191 & ~n13192;
  assign n13194 = ~ a[29]  & ~n13176;
  assign n13195 = ~n13174 & n13177;
  assign n13196 = ~n13194 & ~n13195;
  assign n13197 = n1138 & n3300;
  assign n13198 = n775 & n13197;
  assign n13199 = n288 & n13198;
  assign n13200 = n471 & n13199;
  assign n13201 = n1726 & n13200;
  assign n13202 = n1040 & n13201;
  assign n13203 = ~n752 & n13202;
  assign n13204 = ~n354 & n13203;
  assign n13205 = ~n402 & n13204;
  assign n13206 = ~n505 & n13205;
  assign n13207 = ~n466 & n13206;
  assign n13208 = ~n961 & n13207;
  assign n13209 = ~n332 & n13208;
  assign n13210 = ~n95 & n13209;
  assign n13211 = n621 & n3459;
  assign n13212 = n826 & n13211;
  assign n13213 = ~n713 & n13212;
  assign n13214 = ~n151 & n13213;
  assign n13215 = ~n328 & n13214;
  assign n13216 = ~n417 & n13215;
  assign n13217 = ~n367 & n13216;
  assign n13218 = ~n91 & n13217;
  assign n13219 = ~n132 & n13218;
  assign n13220 = ~n200 & n13219;
  assign n13221 = ~n655 & n13220;
  assign n13222 = n3115 & n5787;
  assign n13223 = n624 & n13222;
  assign n13224 = n494 & n13223;
  assign n13225 = n2987 & n13224;
  assign n13226 = n13221 & n13225;
  assign n13227 = n13210 & n13226;
  assign n13228 = n6707 & n13227;
  assign n13229 = n4232 & n13228;
  assign n13230 = n1254 & n13229;
  assign n13231 = n1531 & n13230;
  assign n13232 = ~n224 & n13231;
  assign n13233 = ~n715 & n13232;
  assign n13234 = ~n568 & n13233;
  assign n13235 = ~n492 & n13234;
  assign n13236 = ~n504 & n13235;
  assign n13237 = ~n453 & n13236;
  assign n13238 = ~n170 & n13237;
  assign n13239 = n13158 & ~n13238;
  assign n13240 = ~n13158 & n13238;
  assign n13241 = n4797 & n12412;
  assign n13242 = n1826 & n13241;
  assign n13243 = n418 & n13242;
  assign n13244 = ~n352 & n13243;
  assign n13245 = ~n144 & n13244;
  assign n13246 = ~n325 & n13245;
  assign n13247 = ~n449 & n13246;
  assign n13248 = ~n146 & ~n713;
  assign n13249 = ~n127 & n13248;
  assign n13250 = n691 & n13249;
  assign n13251 = n6084 & n13250;
  assign n13252 = n6083 & n13251;
  assign n13253 = n1292 & n13252;
  assign n13254 = n3544 & n13253;
  assign n13255 = n285 & n13254;
  assign n13256 = n1825 & n13255;
  assign n13257 = n1366 & n13256;
  assign n13258 = ~n236 & n13257;
  assign n13259 = ~n1306 & n13258;
  assign n13260 = ~n1102 & n13259;
  assign n13261 = ~n287 & n13260;
  assign n13262 = ~n490 & n13261;
  assign n13263 = ~n192 & n13262;
  assign n13264 = ~n246 & n13263;
  assign n13265 = ~n666 & n13264;
  assign n13266 = ~n366 & n590;
  assign n13267 = ~n125 & n13266;
  assign n13268 = ~n428 & n13267;
  assign n13269 = n3645 & n6104;
  assign n13270 = n1557 & n13269;
  assign n13271 = n13268 & n13270;
  assign n13272 = n2772 & n13271;
  assign n13273 = n13265 & n13272;
  assign n13274 = n13247 & n13273;
  assign n13275 = n2090 & n13274;
  assign n13276 = n1330 & n13275;
  assign n13277 = n2406 & n13276;
  assign n13278 = n156 & n13277;
  assign n13279 = n279 & n13278;
  assign n13280 = ~n232 & n13279;
  assign n13281 = ~n327 & n13280;
  assign n13282 = ~n145 & n13281;
  assign n13283 = ~n165 & n13282;
  assign n13284 = ~n12730 & ~n13283;
  assign n13285 = n12730 & n13283;
  assign n13286 = ~n13284 & ~n13285;
  assign n13287 = ~ a[26]  & n13286;
  assign n13288 = ~n13284 & ~n13287;
  assign n13289 = n13238 & ~n13288;
  assign n13290 = n75 & n4477;
  assign n13291 = n3020 & ~n4045;
  assign n13292 = n3023 & ~n3805;
  assign n13293 = n3028 & ~n3964;
  assign n13294 = ~n13292 & ~n13293;
  assign n13295 = ~n13291 & n13294;
  assign n13296 = ~n13290 & n13295;
  assign n13297 = ~n13238 & n13288;
  assign n13298 = ~n13289 & ~n13297;
  assign n13299 = ~n13296 & n13298;
  assign n13300 = ~n13289 & ~n13299;
  assign n13301 = ~n13239 & ~n13300;
  assign n13302 = ~n13240 & n13301;
  assign n13303 = ~n13239 & ~n13302;
  assign n13304 = ~n13196 & ~n13303;
  assign n13305 = n75 & n4715;
  assign n13306 = n3020 & ~n4515;
  assign n13307 = n3023 & ~n4045;
  assign n13308 = n3028 & ~n3877;
  assign n13309 = ~n13307 & ~n13308;
  assign n13310 = ~n13306 & n13309;
  assign n13311 = ~n13305 & n13310;
  assign n13312 = n13196 & n13303;
  assign n13313 = ~n13304 & ~n13312;
  assign n13314 = ~n13311 & n13313;
  assign n13315 = ~n13304 & ~n13314;
  assign n13316 = ~n13193 & ~n13315;
  assign n13317 = n13193 & n13315;
  assign n13318 = ~n13316 & ~n13317;
  assign n13319 = n3542 & ~n4515;
  assign n13320 = n3368 & n4522;
  assign n13321 = ~n13319 & ~n13320;
  assign n13322 =  a[29]  & ~n13321;
  assign n13323 = ~n13321 & ~n13322;
  assign n13324 =  a[29]  & ~n13322;
  assign n13325 = ~n13323 & ~n13324;
  assign n13326 = n75 & n4067;
  assign n13327 = n3020 & ~n3877;
  assign n13328 = n3023 & ~n3964;
  assign n13329 = n3028 & ~n4045;
  assign n13330 = ~n13328 & ~n13329;
  assign n13331 = ~n13327 & n13330;
  assign n13332 = ~n13326 & n13331;
  assign n13333 = ~n13325 & ~n13332;
  assign n13334 = ~n13325 & ~n13333;
  assign n13335 = ~n13332 & ~n13333;
  assign n13336 = ~n13334 & ~n13335;
  assign n13337 = ~n13300 & ~n13302;
  assign n13338 = ~n13240 & n13303;
  assign n13339 = ~n13337 & ~n13338;
  assign n13340 = ~n13336 & ~n13339;
  assign n13341 = ~n13333 & ~n13340;
  assign n13342 = n13311 & ~n13313;
  assign n13343 = ~n13314 & ~n13342;
  assign n13344 = ~n13341 & n13343;
  assign n13345 = ~n13296 & ~n13299;
  assign n13346 = n13298 & ~n13299;
  assign n13347 = ~n13345 & ~n13346;
  assign n13348 = ~ a[26]  & ~n13287;
  assign n13349 = ~n13285 & n13288;
  assign n13350 = ~n13348 & ~n13349;
  assign n13351 = ~n12848 & ~n13350;
  assign n13352 = n75 & n4558;
  assign n13353 = n3020 & ~n3964;
  assign n13354 = n3023 & ~n3456;
  assign n13355 = n3028 & ~n3805;
  assign n13356 = ~n13354 & ~n13355;
  assign n13357 = ~n13353 & n13356;
  assign n13358 = ~n13352 & n13357;
  assign n13359 = n12848 & n13350;
  assign n13360 = ~n13351 & ~n13359;
  assign n13361 = ~n13358 & n13360;
  assign n13362 = ~n13351 & ~n13361;
  assign n13363 = ~n13347 & ~n13362;
  assign n13364 = n13347 & n13362;
  assign n13365 = ~n13363 & ~n13364;
  assign n13366 = n3542 & ~n3877;
  assign n13367 = n3606 & ~n4515;
  assign n13368 = ~n13366 & ~n13367;
  assign n13369 = n3368 & n4609;
  assign n13370 = n13368 & ~n13369;
  assign n13371 =  a[29]  & ~n13370;
  assign n13372 =  a[29]  & ~n13371;
  assign n13373 = ~n13370 & ~n13371;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = n13365 & ~n13374;
  assign n13376 = ~n13363 & ~n13375;
  assign n13377 = ~n13336 & n13339;
  assign n13378 = n13336 & ~n13339;
  assign n13379 = ~n13377 & ~n13378;
  assign n13380 = ~n13376 & ~n13379;
  assign n13381 = n13365 & ~n13375;
  assign n13382 = ~n13374 & ~n13375;
  assign n13383 = ~n13381 & ~n13382;
  assign n13384 = ~n12853 & ~n12856;
  assign n13385 = ~n13358 & ~n13361;
  assign n13386 = n13360 & ~n13361;
  assign n13387 = ~n13385 & ~n13386;
  assign n13388 = ~n13384 & ~n13387;
  assign n13389 = ~n13384 & ~n13388;
  assign n13390 = ~n13387 & ~n13388;
  assign n13391 = ~n13389 & ~n13390;
  assign n13392 = n3457 & ~n4515;
  assign n13393 = n3542 & ~n4045;
  assign n13394 = n3606 & ~n3877;
  assign n13395 = ~n13393 & ~n13394;
  assign n13396 = ~n13392 & n13395;
  assign n13397 = n3368 & n4715;
  assign n13398 = n13396 & ~n13397;
  assign n13399 =  a[29]  & ~n13398;
  assign n13400 =  a[29]  & ~n13399;
  assign n13401 = ~n13398 & ~n13399;
  assign n13402 = ~n13400 & ~n13401;
  assign n13403 = ~n13391 & ~n13402;
  assign n13404 = ~n13388 & ~n13403;
  assign n13405 = ~n13383 & ~n13404;
  assign n13406 = n13383 & n13404;
  assign n13407 = ~n13405 & ~n13406;
  assign n13408 = ~n13391 & ~n13403;
  assign n13409 = ~n13402 & ~n13403;
  assign n13410 = ~n13408 & ~n13409;
  assign n13411 = ~n12877 & ~n12881;
  assign n13412 = ~n13410 & ~n13411;
  assign n13413 = ~n13410 & ~n13412;
  assign n13414 = ~n13411 & ~n13412;
  assign n13415 = ~n13413 & ~n13414;
  assign n13416 = ~n12884 & ~n12887;
  assign n13417 = ~n13415 & ~n13416;
  assign n13418 = ~n13412 & ~n13417;
  assign n13419 = n13407 & ~n13418;
  assign n13420 = ~n13405 & ~n13419;
  assign n13421 = n13376 & n13379;
  assign n13422 = ~n13380 & ~n13421;
  assign n13423 = ~n13420 & n13422;
  assign n13424 = ~n13380 & ~n13423;
  assign n13425 = n13341 & ~n13343;
  assign n13426 = ~n13344 & ~n13425;
  assign n13427 = ~n13424 & n13426;
  assign n13428 = ~n13344 & ~n13427;
  assign n13429 = n13318 & ~n13428;
  assign n13430 = ~n13316 & ~n13429;
  assign n13431 = n13190 & ~n13430;
  assign n13432 = ~n13188 & ~n13431;
  assign n13433 = ~n13109 & ~n13432;
  assign n13434 = ~n13106 & ~n13433;
  assign n13435 = n13059 & ~n13082;
  assign n13436 = ~n13434 & ~n13435;
  assign n13437 = ~n13083 & n13436;
  assign n13438 = ~n13059 & n13437;
  assign n13439 = ~n5407 & ~n5496;
  assign n13440 = ~n4935 & n13439;
  assign n13441 = ~n4938 & n13440;
  assign n13442 = ~n13438 & ~n13441;
  assign n13443 =  a[20]  & ~n13442;
  assign n13444 = ~ a[20]  & n13442;
  assign n13445 = ~n13443 & ~n13444;
  assign n13446 = n336 & n5002;
  assign n13447 = n2595 & n13446;
  assign n13448 = n3435 & n13447;
  assign n13449 = n1894 & n13448;
  assign n13450 = n1245 & n13449;
  assign n13451 = n241 & n13450;
  assign n13452 = n294 & n13451;
  assign n13453 = n1252 & n13452;
  assign n13454 = ~n229 & n13453;
  assign n13455 = ~n232 & n13454;
  assign n13456 = ~n284 & n13455;
  assign n13457 = ~n712 & n13456;
  assign n13458 = ~n562 & n13457;
  assign n13459 = n694 & n3192;
  assign n13460 = n2806 & n13459;
  assign n13461 = n988 & n13460;
  assign n13462 = n805 & n13461;
  assign n13463 = n13458 & n13462;
  assign n13464 = n1708 & n13463;
  assign n13465 = n621 & n13464;
  assign n13466 = n450 & n13465;
  assign n13467 = n869 & n13466;
  assign n13468 = ~n557 & n13467;
  assign n13469 = ~n255 & n13468;
  assign n13470 = ~n252 & n13469;
  assign n13471 = ~n883 & n13470;
  assign n13472 = ~n569 & n13471;
  assign n13473 = ~n771 & n13472;
  assign n13474 = ~n875 & n13473;
  assign n13475 = n12958 & n13474;
  assign n13476 = ~n12958 & ~n13474;
  assign n13477 = ~n13475 & ~n13476;
  assign n13478 = n13445 & n13477;
  assign n13479 = ~n13445 & ~n13477;
  assign n13480 = ~n13478 & ~n13479;
  assign n13481 = ~n13009 & n13480;
  assign n13482 = n13009 & ~n13480;
  assign n13483 = ~n13481 & ~n13482;
  assign n13484 = ~n12902 & n13483;
  assign n13485 = ~n13481 & ~n13484;
  assign n13486 = ~n13476 & ~n13478;
  assign n13487 = n13031 & ~n13486;
  assign n13488 = ~n13031 & n13486;
  assign n13489 = ~n13487 & ~n13488;
  assign n13490 = n13415 & n13416;
  assign n13491 = ~n13417 & ~n13490;
  assign n13492 = n3020 & n13491;
  assign n13493 = n3028 & n12889;
  assign n13494 = n3023 & n12769;
  assign n13495 = ~n12891 & ~n12893;
  assign n13496 = n12889 & n13491;
  assign n13497 = ~n12889 & ~n13491;
  assign n13498 = ~n13495 & ~n13497;
  assign n13499 = ~n13496 & n13498;
  assign n13500 = ~n13495 & ~n13499;
  assign n13501 = ~n13496 & ~n13499;
  assign n13502 = ~n13497 & n13501;
  assign n13503 = ~n13500 & ~n13502;
  assign n13504 = n75 & ~n13503;
  assign n13505 = ~n13494 & ~n13504;
  assign n13506 = ~n13493 & n13505;
  assign n13507 = ~n13492 & n13506;
  assign n13508 = n13489 & ~n13507;
  assign n13509 = ~n13489 & n13507;
  assign n13510 = ~n13508 & ~n13509;
  assign n13511 = ~n13485 & n13510;
  assign n13512 = n13485 & ~n13510;
  assign n13513 = ~n13511 & ~n13512;
  assign n13514 = n13424 & ~n13426;
  assign n13515 = ~n13427 & ~n13514;
  assign n13516 = n3457 & n13515;
  assign n13517 = ~n13407 & n13418;
  assign n13518 = ~n13419 & ~n13517;
  assign n13519 = n3542 & n13518;
  assign n13520 = n13420 & ~n13422;
  assign n13521 = ~n13423 & ~n13520;
  assign n13522 = n3606 & n13521;
  assign n13523 = ~n13519 & ~n13522;
  assign n13524 = ~n13516 & n13523;
  assign n13525 = ~n3368 & n13524;
  assign n13526 = n13518 & n13521;
  assign n13527 = n13491 & n13518;
  assign n13528 = ~n13491 & ~n13518;
  assign n13529 = ~n13527 & ~n13528;
  assign n13530 = ~n13501 & n13529;
  assign n13531 = ~n13527 & ~n13530;
  assign n13532 = ~n13518 & ~n13521;
  assign n13533 = ~n13531 & ~n13532;
  assign n13534 = ~n13526 & n13533;
  assign n13535 = ~n13526 & ~n13534;
  assign n13536 = ~n13515 & ~n13521;
  assign n13537 = n13515 & n13521;
  assign n13538 = ~n13536 & ~n13537;
  assign n13539 = ~n13535 & n13538;
  assign n13540 = n13535 & ~n13538;
  assign n13541 = ~n13539 & ~n13540;
  assign n13542 = n13524 & ~n13541;
  assign n13543 = ~n13525 & ~n13542;
  assign n13544 =  a[29]  & ~n13543;
  assign n13545 = ~ a[29]  & n13543;
  assign n13546 = ~n13544 & ~n13545;
  assign n13547 = n13513 & ~n13546;
  assign n13548 = ~n13511 & ~n13547;
  assign n13549 = ~n13487 & ~n13508;
  assign n13550 = n3792 & n4788;
  assign n13551 = n989 & n13550;
  assign n13552 = n2371 & n13551;
  assign n13553 = n3544 & n13552;
  assign n13554 = n285 & n13553;
  assign n13555 = ~n398 & n13554;
  assign n13556 = ~n1062 & n13555;
  assign n13557 = ~n619 & n13556;
  assign n13558 = ~n470 & n13557;
  assign n13559 = ~n271 & n13558;
  assign n13560 = ~n125 & n13559;
  assign n13561 = n3549 & n5734;
  assign n13562 = n12390 & n13561;
  assign n13563 = n3389 & n13562;
  assign n13564 = n12939 & n13563;
  assign n13565 = n13560 & n13564;
  assign n13566 = n4293 & n13565;
  assign n13567 = n2021 & n13566;
  assign n13568 = n896 & n13567;
  assign n13569 = n3886 & n13568;
  assign n13570 = ~n847 & n13569;
  assign n13571 = ~n175 & n13570;
  assign n13572 = ~n286 & n13571;
  assign n13573 = ~n563 & n13572;
  assign n13574 = ~n368 & n13573;
  assign n13575 = ~n13031 & n13574;
  assign n13576 = n13031 & ~n13574;
  assign n13577 = ~n13549 & ~n13576;
  assign n13578 = ~n13575 & n13577;
  assign n13579 = ~n13549 & ~n13578;
  assign n13580 = ~n13575 & ~n13578;
  assign n13581 = ~n13576 & n13580;
  assign n13582 = ~n13579 & ~n13581;
  assign n13583 = n13501 & ~n13529;
  assign n13584 = ~n13530 & ~n13583;
  assign n13585 = n75 & n13584;
  assign n13586 = n3020 & n13518;
  assign n13587 = n3023 & n12889;
  assign n13588 = n3028 & n13491;
  assign n13589 = ~n13587 & ~n13588;
  assign n13590 = ~n13586 & n13589;
  assign n13591 = ~n13585 & n13590;
  assign n13592 = ~n13582 & ~n13591;
  assign n13593 = ~n13582 & ~n13592;
  assign n13594 = ~n13591 & ~n13592;
  assign n13595 = ~n13593 & ~n13594;
  assign n13596 = ~n13318 & n13428;
  assign n13597 = ~n13429 & ~n13596;
  assign n13598 = n3457 & n13597;
  assign n13599 = n3542 & n13521;
  assign n13600 = n3606 & n13515;
  assign n13601 = ~n13599 & ~n13600;
  assign n13602 = ~n13598 & n13601;
  assign n13603 = ~n3368 & n13602;
  assign n13604 = ~n13537 & ~n13539;
  assign n13605 = n13515 & n13597;
  assign n13606 = ~n13515 & ~n13597;
  assign n13607 = ~n13604 & ~n13606;
  assign n13608 = ~n13605 & n13607;
  assign n13609 = ~n13604 & ~n13608;
  assign n13610 = ~n13605 & ~n13608;
  assign n13611 = ~n13606 & n13610;
  assign n13612 = ~n13609 & ~n13611;
  assign n13613 = n13602 & n13612;
  assign n13614 = ~n13603 & ~n13613;
  assign n13615 =  a[29]  & ~n13614;
  assign n13616 = ~ a[29]  & n13614;
  assign n13617 = ~n13615 & ~n13616;
  assign n13618 = ~n13595 & ~n13617;
  assign n13619 = n13595 & n13617;
  assign n13620 = ~n13618 & ~n13619;
  assign n13621 = ~n13548 & n13620;
  assign n13622 = n13548 & ~n13620;
  assign n13623 = ~n13621 & ~n13622;
  assign n13624 = ~n13434 & ~n13437;
  assign n13625 = ~n13435 & ~n13437;
  assign n13626 = ~n13083 & n13625;
  assign n13627 = ~n13624 & ~n13626;
  assign n13628 = n3884 & ~n13627;
  assign n13629 = ~n13190 & n13430;
  assign n13630 = ~n13431 & ~n13629;
  assign n13631 = n3967 & n13630;
  assign n13632 = n13109 & n13432;
  assign n13633 = ~n13433 & ~n13632;
  assign n13634 = n4046 & n13633;
  assign n13635 = ~n13631 & ~n13634;
  assign n13636 = ~n13628 & n13635;
  assign n13637 = n13630 & n13633;
  assign n13638 = n13597 & n13630;
  assign n13639 = ~n13597 & ~n13630;
  assign n13640 = ~n13638 & ~n13639;
  assign n13641 = ~n13610 & n13640;
  assign n13642 = ~n13638 & ~n13641;
  assign n13643 = ~n13630 & ~n13633;
  assign n13644 = ~n13637 & ~n13643;
  assign n13645 = ~n13642 & n13644;
  assign n13646 = ~n13637 & ~n13645;
  assign n13647 = ~n13627 & n13633;
  assign n13648 = n13627 & ~n13633;
  assign n13649 = ~n13646 & ~n13648;
  assign n13650 = ~n13647 & n13649;
  assign n13651 = ~n13646 & ~n13650;
  assign n13652 = ~n13647 & ~n13650;
  assign n13653 = ~n13648 & n13652;
  assign n13654 = ~n13651 & ~n13653;
  assign n13655 = n4050 & ~n13654;
  assign n13656 = n13636 & ~n13655;
  assign n13657 =  a[26]  & ~n13656;
  assign n13658 =  a[26]  & ~n13657;
  assign n13659 = ~n13656 & ~n13657;
  assign n13660 = ~n13658 & ~n13659;
  assign n13661 = n13623 & ~n13660;
  assign n13662 = n13623 & ~n13661;
  assign n13663 = ~n13660 & ~n13661;
  assign n13664 = ~n13662 & ~n13663;
  assign n13665 = n13483 & ~n13484;
  assign n13666 = ~n12902 & ~n13484;
  assign n13667 = ~n13665 & ~n13666;
  assign n13668 = ~n13006 & ~n13008;
  assign n13669 = ~n12997 & n13009;
  assign n13670 = ~n13668 & ~n13669;
  assign n13671 = ~n330 & ~n352;
  assign n13672 = ~n1072 & n2809;
  assign n13673 = ~n847 & n13672;
  assign n13674 = ~n557 & n13673;
  assign n13675 = ~n417 & n13674;
  assign n13676 = ~n568 & n13675;
  assign n13677 = ~n205 & n13676;
  assign n13678 = n1437 & n2220;
  assign n13679 = n2487 & n13678;
  assign n13680 = n2345 & n13679;
  assign n13681 = n13677 & n13680;
  assign n13682 = n772 & n13681;
  assign n13683 = n3108 & n13682;
  assign n13684 = n5264 & n13683;
  assign n13685 = n4786 & n13684;
  assign n13686 = n1824 & n13685;
  assign n13687 = n2583 & n13686;
  assign n13688 = n2466 & n13687;
  assign n13689 = ~n189 & n13688;
  assign n13690 = n13671 & n13689;
  assign n13691 = ~n656 & n13690;
  assign n13692 = ~n492 & n13691;
  assign n13693 = ~n201 & n13692;
  assign n13694 = ~n470 & n13693;
  assign n13695 = ~n86 & n13694;
  assign n13696 = ~n656 & ~n809;
  assign n13697 = ~n145 & n13696;
  assign n13698 = ~n489 & n13697;
  assign n13699 = n421 & ~n639;
  assign n13700 = ~n592 & n13699;
  assign n13701 = n2753 & n13700;
  assign n13702 = n6672 & n13701;
  assign n13703 = n13138 & n13702;
  assign n13704 = n13698 & n13703;
  assign n13705 = n12919 & n13704;
  assign n13706 = n4815 & n13705;
  assign n13707 = n2605 & n13706;
  assign n13708 = n1575 & n13707;
  assign n13709 = n2406 & n13708;
  assign n13710 = n202 & n13709;
  assign n13711 = n1380 & n13710;
  assign n13712 = ~n136 & n13711;
  assign n13713 = ~n327 & n13712;
  assign n13714 = ~n393 & n13713;
  assign n13715 = ~n270 & n13714;
  assign n13716 = ~n13695 & ~n13715;
  assign n13717 = ~n5939 & ~n6233;
  assign n13718 = ~n5663 & n13717;
  assign n13719 = ~n5666 & n13718;
  assign n13720 = ~n13438 & ~n13719;
  assign n13721 =  a[17]  & ~n13720;
  assign n13722 = ~ a[17]  & n13720;
  assign n13723 = ~n13721 & ~n13722;
  assign n13724 = n13695 & n13715;
  assign n13725 = ~n13716 & ~n13724;
  assign n13726 = n13723 & n13725;
  assign n13727 = ~n13716 & ~n13726;
  assign n13728 = n12958 & ~n13727;
  assign n13729 = ~n12958 & n13727;
  assign n13730 = ~n13728 & ~n13729;
  assign n13731 = n3020 & n12502;
  assign n13732 = n3028 & n12370;
  assign n13733 = n3023 & n12505;
  assign n13734 = ~n12680 & ~n12683;
  assign n13735 = ~n12681 & n12684;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = n75 & ~n13736;
  assign n13738 = ~n13733 & ~n13737;
  assign n13739 = ~n13732 & n13738;
  assign n13740 = ~n13731 & n13739;
  assign n13741 = n13730 & ~n13740;
  assign n13742 = ~n13728 & ~n13741;
  assign n13743 = ~n13670 & ~n13742;
  assign n13744 = n13670 & n13742;
  assign n13745 = ~n13743 & ~n13744;
  assign n13746 = ~n12676 & ~n12679;
  assign n13747 = ~n12677 & n12680;
  assign n13748 = ~n13746 & ~n13747;
  assign n13749 = n75 & ~n13748;
  assign n13750 = n3020 & n12370;
  assign n13751 = n3023 & n12508;
  assign n13752 = n3028 & n12505;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = ~n13750 & n13753;
  assign n13755 = ~n13749 & n13754;
  assign n13756 = ~n13723 & ~n13725;
  assign n13757 = ~n13726 & ~n13756;
  assign n13758 = ~n13755 & n13757;
  assign n13759 = n1253 & n2739;
  assign n13760 = n2090 & n13759;
  assign n13761 = n238 & n13760;
  assign n13762 = ~n427 & n13761;
  assign n13763 = ~n335 & n13762;
  assign n13764 = ~n280 & n13763;
  assign n13765 = ~n239 & n13764;
  assign n13766 = ~n460 & n13765;
  assign n13767 = ~n657 & n13766;
  assign n13768 = ~n86 & n13767;
  assign n13769 = ~n617 & ~n1306;
  assign n13770 = ~n752 & n13769;
  assign n13771 = ~n602 & n13770;
  assign n13772 = ~n286 & n13771;
  assign n13773 = ~n532 & n13772;
  assign n13774 = ~n130 & ~n144;
  assign n13775 = n3160 & n13774;
  assign n13776 = n13773 & n13775;
  assign n13777 = n4325 & n13776;
  assign n13778 = n6020 & n13777;
  assign n13779 = n1366 & n13778;
  assign n13780 = ~n667 & n13779;
  assign n13781 = ~n232 & n13780;
  assign n13782 = ~n495 & n13781;
  assign n13783 = ~n435 & n13782;
  assign n13784 = ~n248 & n13783;
  assign n13785 = ~n91 & n13784;
  assign n13786 = ~n272 & n13785;
  assign n13787 = ~n886 & n13786;
  assign n13788 = n2683 & n13787;
  assign n13789 = ~n168 & n13788;
  assign n13790 = n1308 & n13789;
  assign n13791 = n1942 & n13790;
  assign n13792 = n5791 & n13791;
  assign n13793 = n2796 & n13792;
  assign n13794 = n13768 & n13793;
  assign n13795 = n1575 & n13794;
  assign n13796 = n2484 & n13795;
  assign n13797 = n159 & n13796;
  assign n13798 = n1161 & n13797;
  assign n13799 = ~n229 & n13798;
  assign n13800 = ~n329 & n13799;
  assign n13801 = ~n353 & n13800;
  assign n13802 = ~n639 & n13801;
  assign n13803 = ~n567 & n13802;
  assign n13804 = ~n712 & n13803;
  assign n13805 = ~n304 & n13804;
  assign n13806 = n13695 & ~n13805;
  assign n13807 = ~n136 & n5082;
  assign n13808 = ~n884 & n13807;
  assign n13809 = n5271 & n13808;
  assign n13810 = n3041 & n13809;
  assign n13811 = n2716 & n13810;
  assign n13812 = n3489 & n13811;
  assign n13813 = n4367 & n13812;
  assign n13814 = n1080 & n13813;
  assign n13815 = ~n518 & n13814;
  assign n13816 = ~n602 & n13815;
  assign n13817 = ~n146 & n13816;
  assign n13818 = n888 & n13817;
  assign n13819 = ~n673 & n13818;
  assign n13820 = ~n564 & n13819;
  assign n13821 = ~n125 & n13820;
  assign n13822 = n423 & n1366;
  assign n13823 = ~n151 & n13822;
  assign n13824 = ~n537 & n13823;
  assign n13825 = ~n375 & n13824;
  assign n13826 = ~n222 & n13825;
  assign n13827 = n773 & n1528;
  assign n13828 = n1346 & n13827;
  assign n13829 = n4298 & n13828;
  assign n13830 = n3068 & n13829;
  assign n13831 = n434 & n13830;
  assign n13832 = n13826 & n13831;
  assign n13833 = n1814 & n13832;
  assign n13834 = n6514 & n13833;
  assign n13835 = n774 & n13834;
  assign n13836 = n1838 & n13835;
  assign n13837 = ~n232 & n13836;
  assign n13838 = ~n637 & n13837;
  assign n13839 = ~n228 & n13838;
  assign n13840 = ~n302 & n13839;
  assign n13841 = ~n298 & n13840;
  assign n13842 = ~n295 & n13841;
  assign n13843 = ~n127 & n13842;
  assign n13844 = ~n13821 & ~n13843;
  assign n13845 = ~n6951 & ~n7101;
  assign n13846 = ~n6402 & n13845;
  assign n13847 = ~n6397 & n13846;
  assign n13848 = ~n13438 & ~n13847;
  assign n13849 =  a[14]  & ~n13848;
  assign n13850 = ~ a[14]  & n13848;
  assign n13851 = ~n13849 & ~n13850;
  assign n13852 = n13821 & n13843;
  assign n13853 = ~n13844 & ~n13852;
  assign n13854 = n13851 & n13853;
  assign n13855 = ~n13844 & ~n13854;
  assign n13856 = n13805 & ~n13855;
  assign n13857 = ~n13805 & n13855;
  assign n13858 = ~n13856 & ~n13857;
  assign n13859 = n3020 & n12508;
  assign n13860 = n3028 & n12513;
  assign n13861 = n3023 & n12511;
  assign n13862 = n12667 & ~n12670;
  assign n13863 = ~n12671 & ~n13862;
  assign n13864 = n75 & n13863;
  assign n13865 = ~n13861 & ~n13864;
  assign n13866 = ~n13860 & n13865;
  assign n13867 = ~n13859 & n13866;
  assign n13868 = n13858 & ~n13867;
  assign n13869 = ~n13856 & ~n13868;
  assign n13870 = ~n13695 & n13805;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = ~n13806 & n13871;
  assign n13873 = ~n13806 & ~n13872;
  assign n13874 = n13757 & ~n13758;
  assign n13875 = ~n13755 & ~n13758;
  assign n13876 = ~n13874 & ~n13875;
  assign n13877 = ~n13873 & ~n13876;
  assign n13878 = ~n13758 & ~n13877;
  assign n13879 = ~n13730 & n13740;
  assign n13880 = ~n13741 & ~n13879;
  assign n13881 = ~n13878 & n13880;
  assign n13882 = n13878 & ~n13880;
  assign n13883 = ~n13881 & ~n13882;
  assign n13884 = n3457 & n13491;
  assign n13885 = n3542 & n12769;
  assign n13886 = n3606 & n12889;
  assign n13887 = ~n13885 & ~n13886;
  assign n13888 = ~n13884 & n13887;
  assign n13889 = ~n3368 & n13888;
  assign n13890 = n13503 & n13888;
  assign n13891 = ~n13889 & ~n13890;
  assign n13892 =  a[29]  & ~n13891;
  assign n13893 = ~ a[29]  & n13891;
  assign n13894 = ~n13892 & ~n13893;
  assign n13895 = n13883 & ~n13894;
  assign n13896 = ~n13881 & ~n13895;
  assign n13897 = n13745 & ~n13896;
  assign n13898 = ~n13743 & ~n13897;
  assign n13899 = ~n13667 & ~n13898;
  assign n13900 = n13667 & n13898;
  assign n13901 = ~n13899 & ~n13900;
  assign n13902 = n3457 & n13521;
  assign n13903 = n3542 & n13491;
  assign n13904 = n3606 & n13518;
  assign n13905 = ~n13903 & ~n13904;
  assign n13906 = ~n13902 & n13905;
  assign n13907 = ~n13531 & ~n13534;
  assign n13908 = ~n13532 & n13535;
  assign n13909 = ~n13907 & ~n13908;
  assign n13910 = n3368 & ~n13909;
  assign n13911 = n13906 & ~n13910;
  assign n13912 =  a[29]  & ~n13911;
  assign n13913 =  a[29]  & ~n13912;
  assign n13914 = ~n13911 & ~n13912;
  assign n13915 = ~n13913 & ~n13914;
  assign n13916 = n13901 & ~n13915;
  assign n13917 = ~n13899 & ~n13916;
  assign n13918 = ~n13513 & n13546;
  assign n13919 = ~n13547 & ~n13918;
  assign n13920 = ~n13917 & n13919;
  assign n13921 = n13917 & ~n13919;
  assign n13922 = ~n13920 & ~n13921;
  assign n13923 = n3884 & n13633;
  assign n13924 = n3967 & n13597;
  assign n13925 = n4046 & n13630;
  assign n13926 = ~n13924 & ~n13925;
  assign n13927 = ~n13923 & n13926;
  assign n13928 = n13642 & ~n13644;
  assign n13929 = ~n13645 & ~n13928;
  assign n13930 = n4050 & n13929;
  assign n13931 = n13927 & ~n13930;
  assign n13932 =  a[26]  & ~n13931;
  assign n13933 =  a[26]  & ~n13932;
  assign n13934 = ~n13931 & ~n13932;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = n13922 & ~n13935;
  assign n13937 = ~n13920 & ~n13936;
  assign n13938 = ~n4604 & ~n4694;
  assign n13939 = ~n13438 & ~n13938;
  assign n13940 = n13059 & n13625;
  assign n13941 = ~n13438 & ~n13940;
  assign n13942 = n4533 & n13941;
  assign n13943 = ~n13939 & ~n13942;
  assign n13944 = ~n4536 & n13943;
  assign n13945 = ~n13627 & n13941;
  assign n13946 = n13627 & ~n13941;
  assign n13947 = ~n13945 & ~n13946;
  assign n13948 = ~n13652 & n13947;
  assign n13949 = ~n13945 & ~n13948;
  assign n13950 = n13940 & ~n13949;
  assign n13951 = ~n13941 & ~n13950;
  assign n13952 = n13943 & n13951;
  assign n13953 = ~n13944 & ~n13952;
  assign n13954 =  a[23]  & ~n13953;
  assign n13955 = ~ a[23]  & n13953;
  assign n13956 = ~n13954 & ~n13955;
  assign n13957 = ~n13937 & ~n13956;
  assign n13958 = n13937 & n13956;
  assign n13959 = ~n13957 & ~n13958;
  assign n13960 = ~n13664 & n13959;
  assign n13961 = ~n13664 & ~n13960;
  assign n13962 = n13959 & ~n13960;
  assign n13963 = ~n13961 & ~n13962;
  assign n13964 = n13922 & ~n13936;
  assign n13965 = ~n13935 & ~n13936;
  assign n13966 = ~n13964 & ~n13965;
  assign n13967 = n13901 & ~n13916;
  assign n13968 = ~n13915 & ~n13916;
  assign n13969 = ~n13967 & ~n13968;
  assign n13970 = n3884 & n13630;
  assign n13971 = n3967 & n13515;
  assign n13972 = n4046 & n13597;
  assign n13973 = ~n13971 & ~n13972;
  assign n13974 = ~n13970 & n13973;
  assign n13975 = n13610 & ~n13640;
  assign n13976 = ~n13641 & ~n13975;
  assign n13977 = n4050 & n13976;
  assign n13978 = n13974 & ~n13977;
  assign n13979 =  a[26]  & ~n13978;
  assign n13980 =  a[26]  & ~n13979;
  assign n13981 = ~n13978 & ~n13979;
  assign n13982 = ~n13980 & ~n13981;
  assign n13983 = ~n13969 & ~n13982;
  assign n13984 = ~n13969 & ~n13983;
  assign n13985 = ~n13982 & ~n13983;
  assign n13986 = ~n13984 & ~n13985;
  assign n13987 = ~n13745 & n13896;
  assign n13988 = ~n13897 & ~n13987;
  assign n13989 = n3457 & n13518;
  assign n13990 = n3542 & n12889;
  assign n13991 = n3606 & n13491;
  assign n13992 = ~n13990 & ~n13991;
  assign n13993 = ~n13989 & n13992;
  assign n13994 = n3368 & n13584;
  assign n13995 = n13993 & ~n13994;
  assign n13996 =  a[29]  & ~n13995;
  assign n13997 =  a[29]  & ~n13996;
  assign n13998 = ~n13995 & ~n13996;
  assign n13999 = ~n13997 & ~n13998;
  assign n14000 = n13988 & ~n13999;
  assign n14001 = n13988 & ~n14000;
  assign n14002 = ~n13999 & ~n14000;
  assign n14003 = ~n14001 & ~n14002;
  assign n14004 = n3884 & n13597;
  assign n14005 = n3967 & n13521;
  assign n14006 = n4046 & n13515;
  assign n14007 = ~n14005 & ~n14006;
  assign n14008 = ~n14004 & n14007;
  assign n14009 = n4050 & ~n13612;
  assign n14010 = n14008 & ~n14009;
  assign n14011 =  a[26]  & ~n14010;
  assign n14012 =  a[26]  & ~n14011;
  assign n14013 = ~n14010 & ~n14011;
  assign n14014 = ~n14012 & ~n14013;
  assign n14015 = ~n14003 & ~n14014;
  assign n14016 = ~n14000 & ~n14015;
  assign n14017 = ~n13986 & ~n14016;
  assign n14018 = ~n13983 & ~n14017;
  assign n14019 = ~n13966 & ~n14018;
  assign n14020 = n13966 & n14018;
  assign n14021 = ~n14019 & ~n14020;
  assign n14022 = n4694 & ~n13438;
  assign n14023 = n4533 & ~n13627;
  assign n14024 = n4604 & n13941;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = ~n14022 & n14025;
  assign n14027 = ~n13940 & n13949;
  assign n14028 = ~n13950 & ~n14027;
  assign n14029 = n4536 & n14028;
  assign n14030 = n14026 & ~n14029;
  assign n14031 =  a[23]  & ~n14030;
  assign n14032 =  a[23]  & ~n14031;
  assign n14033 = ~n14030 & ~n14031;
  assign n14034 = ~n14032 & ~n14033;
  assign n14035 = n14021 & ~n14034;
  assign n14036 = ~n14019 & ~n14035;
  assign n14037 = ~n13963 & ~n14036;
  assign n14038 = n13963 & n14036;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = n14021 & ~n14035;
  assign n14041 = ~n14034 & ~n14035;
  assign n14042 = ~n14040 & ~n14041;
  assign n14043 = ~n14003 & ~n14015;
  assign n14044 = ~n14014 & ~n14015;
  assign n14045 = ~n14043 & ~n14044;
  assign n14046 = ~n13869 & ~n13872;
  assign n14047 = ~n13870 & n13873;
  assign n14048 = ~n14046 & ~n14047;
  assign n14049 = ~n12672 & ~n12675;
  assign n14050 = ~n12673 & n12676;
  assign n14051 = ~n14049 & ~n14050;
  assign n14052 = n75 & ~n14051;
  assign n14053 = n3020 & n12505;
  assign n14054 = n3023 & n12513;
  assign n14055 = n3028 & n12508;
  assign n14056 = ~n14054 & ~n14055;
  assign n14057 = ~n14053 & n14056;
  assign n14058 = ~n14052 & n14057;
  assign n14059 = ~n14048 & ~n14058;
  assign n14060 = ~n14048 & ~n14059;
  assign n14061 = ~n14058 & ~n14059;
  assign n14062 = ~n14060 & ~n14061;
  assign n14063 = n3457 & n12769;
  assign n14064 = n3542 & n12370;
  assign n14065 = n3606 & n12502;
  assign n14066 = ~n14064 & ~n14065;
  assign n14067 = ~n14063 & n14066;
  assign n14068 = ~n3368 & n14067;
  assign n14069 = ~n12999 & n14067;
  assign n14070 = ~n14068 & ~n14069;
  assign n14071 =  a[29]  & ~n14070;
  assign n14072 = ~ a[29]  & n14070;
  assign n14073 = ~n14071 & ~n14072;
  assign n14074 = ~n14062 & ~n14073;
  assign n14075 = ~n14059 & ~n14074;
  assign n14076 = ~n13876 & ~n13877;
  assign n14077 = ~n13873 & ~n13877;
  assign n14078 = ~n14076 & ~n14077;
  assign n14079 = ~n14075 & ~n14078;
  assign n14080 = ~n14075 & ~n14079;
  assign n14081 = ~n14078 & ~n14079;
  assign n14082 = ~n14080 & ~n14081;
  assign n14083 = n3457 & n12889;
  assign n14084 = n3542 & n12502;
  assign n14085 = n3606 & n12769;
  assign n14086 = ~n14084 & ~n14085;
  assign n14087 = ~n14083 & n14086;
  assign n14088 = n3368 & n12895;
  assign n14089 = n14087 & ~n14088;
  assign n14090 =  a[29]  & ~n14089;
  assign n14091 =  a[29]  & ~n14090;
  assign n14092 = ~n14089 & ~n14090;
  assign n14093 = ~n14091 & ~n14092;
  assign n14094 = ~n14082 & ~n14093;
  assign n14095 = ~n14079 & ~n14094;
  assign n14096 = ~n13883 & n13894;
  assign n14097 = ~n13895 & ~n14096;
  assign n14098 = ~n14095 & n14097;
  assign n14099 = n14095 & ~n14097;
  assign n14100 = ~n14098 & ~n14099;
  assign n14101 = n3884 & n13515;
  assign n14102 = n3967 & n13518;
  assign n14103 = n4046 & n13521;
  assign n14104 = ~n14102 & ~n14103;
  assign n14105 = ~n14101 & n14104;
  assign n14106 = n4050 & n13541;
  assign n14107 = n14105 & ~n14106;
  assign n14108 =  a[26]  & ~n14107;
  assign n14109 =  a[26]  & ~n14108;
  assign n14110 = ~n14107 & ~n14108;
  assign n14111 = ~n14109 & ~n14110;
  assign n14112 = n14100 & ~n14111;
  assign n14113 = ~n14098 & ~n14112;
  assign n14114 = ~n14045 & ~n14113;
  assign n14115 = n14045 & n14113;
  assign n14116 = ~n14114 & ~n14115;
  assign n14117 = n4694 & ~n13627;
  assign n14118 = n4533 & n13630;
  assign n14119 = n4604 & n13633;
  assign n14120 = ~n14118 & ~n14119;
  assign n14121 = ~n14117 & n14120;
  assign n14122 = n4536 & ~n13654;
  assign n14123 = n14121 & ~n14122;
  assign n14124 =  a[23]  & ~n14123;
  assign n14125 =  a[23]  & ~n14124;
  assign n14126 = ~n14123 & ~n14124;
  assign n14127 = ~n14125 & ~n14126;
  assign n14128 = n14116 & ~n14127;
  assign n14129 = ~n14114 & ~n14128;
  assign n14130 = n4694 & n13941;
  assign n14131 = n4533 & n13633;
  assign n14132 = n4604 & ~n13627;
  assign n14133 = ~n14131 & ~n14132;
  assign n14134 = ~n14130 & n14133;
  assign n14135 = n13652 & ~n13947;
  assign n14136 = ~n13948 & ~n14135;
  assign n14137 = n4536 & n14136;
  assign n14138 = n14134 & ~n14137;
  assign n14139 =  a[23]  & ~n14138;
  assign n14140 =  a[23]  & ~n14139;
  assign n14141 = ~n14138 & ~n14139;
  assign n14142 = ~n14140 & ~n14141;
  assign n14143 = ~n14129 & ~n14142;
  assign n14144 = n13986 & n14016;
  assign n14145 = ~n14017 & ~n14144;
  assign n14146 = ~n14129 & ~n14143;
  assign n14147 = ~n14142 & ~n14143;
  assign n14148 = ~n14146 & ~n14147;
  assign n14149 = n14145 & ~n14148;
  assign n14150 = ~n14143 & ~n14149;
  assign n14151 = ~n14042 & ~n14150;
  assign n14152 = ~n14042 & ~n14151;
  assign n14153 = ~n14150 & ~n14151;
  assign n14154 = ~n14152 & ~n14153;
  assign n14155 = n14100 & ~n14112;
  assign n14156 = ~n14111 & ~n14112;
  assign n14157 = ~n14155 & ~n14156;
  assign n14158 = ~n14082 & ~n14094;
  assign n14159 = ~n14093 & ~n14094;
  assign n14160 = ~n14158 & ~n14159;
  assign n14161 = n3884 & n13521;
  assign n14162 = n3967 & n13491;
  assign n14163 = n4046 & n13518;
  assign n14164 = ~n14162 & ~n14163;
  assign n14165 = ~n14161 & n14164;
  assign n14166 = n4050 & ~n13909;
  assign n14167 = n14165 & ~n14166;
  assign n14168 =  a[26]  & ~n14167;
  assign n14169 =  a[26]  & ~n14168;
  assign n14170 = ~n14167 & ~n14168;
  assign n14171 = ~n14169 & ~n14170;
  assign n14172 = ~n14160 & ~n14171;
  assign n14173 = ~n14160 & ~n14172;
  assign n14174 = ~n14171 & ~n14172;
  assign n14175 = ~n14173 & ~n14174;
  assign n14176 = n12663 & ~n12665;
  assign n14177 = ~n12666 & ~n14176;
  assign n14178 = n75 & n14177;
  assign n14179 = n3020 & n12513;
  assign n14180 = n3023 & n12516;
  assign n14181 = n3028 & n12511;
  assign n14182 = ~n14180 & ~n14181;
  assign n14183 = ~n14179 & n14182;
  assign n14184 = ~n14178 & n14183;
  assign n14185 = ~n142 & ~n506;
  assign n14186 = ~n422 & n14185;
  assign n14187 = ~n603 & n14186;
  assign n14188 = ~n130 & n14187;
  assign n14189 = ~n332 & n14188;
  assign n14190 = n1109 & n3523;
  assign n14191 = n5777 & n14190;
  assign n14192 = n14189 & n14191;
  assign n14193 = n2022 & n14192;
  assign n14194 = n622 & n14193;
  assign n14195 = n874 & n14194;
  assign n14196 = n774 & n14195;
  assign n14197 = n872 & n14196;
  assign n14198 = n356 & n14197;
  assign n14199 = ~n1306 & n14198;
  assign n14200 = ~n403 & n14199;
  assign n14201 = ~n161 & n14200;
  assign n14202 = ~n655 & n14201;
  assign n14203 = n642 & n3165;
  assign n14204 = n2390 & n14203;
  assign n14205 = n989 & n14204;
  assign n14206 = n1782 & n14205;
  assign n14207 = ~n1011 & n14206;
  assign n14208 = ~n847 & n14207;
  assign n14209 = ~n331 & n14208;
  assign n14210 = ~n132 & n14209;
  assign n14211 = n529 & n14210;
  assign n14212 = n3681 & n14211;
  assign n14213 = n2296 & n14212;
  assign n14214 = n14202 & n14213;
  assign n14215 = n1046 & n14214;
  assign n14216 = n450 & n14215;
  assign n14217 = n937 & n14216;
  assign n14218 = n2088 & n14217;
  assign n14219 = n4101 & n14218;
  assign n14220 = n1522 & n14219;
  assign n14221 = ~n136 & n14220;
  assign n14222 = ~n1062 & n14221;
  assign n14223 = ~n302 & n14222;
  assign n14224 = ~n192 & n14223;
  assign n14225 = ~n430 & n14224;
  assign n14226 = ~n201 & n14225;
  assign n14227 = ~n657 & n14226;
  assign n14228 = ~n158 & n14227;
  assign n14229 = n13821 & ~n14228;
  assign n14230 = ~n13821 & n14228;
  assign n14231 = ~n12659 & ~n12662;
  assign n14232 = ~n12660 & n12663;
  assign n14233 = ~n14231 & ~n14232;
  assign n14234 = n75 & ~n14233;
  assign n14235 = n3020 & n12511;
  assign n14236 = n3023 & n12519;
  assign n14237 = n3028 & n12516;
  assign n14238 = ~n14236 & ~n14237;
  assign n14239 = ~n14235 & n14238;
  assign n14240 = ~n14234 & n14239;
  assign n14241 = ~n14229 & ~n14240;
  assign n14242 = ~n14230 & n14241;
  assign n14243 = ~n14229 & ~n14242;
  assign n14244 = ~n13851 & ~n13853;
  assign n14245 = ~n13854 & ~n14244;
  assign n14246 = ~n14243 & n14245;
  assign n14247 = n14243 & ~n14245;
  assign n14248 = ~n14246 & ~n14247;
  assign n14249 = ~n14184 & n14248;
  assign n14250 = ~n14246 & ~n14249;
  assign n14251 = ~n13858 & n13867;
  assign n14252 = ~n13868 & ~n14251;
  assign n14253 = ~n14250 & n14252;
  assign n14254 = n14250 & ~n14252;
  assign n14255 = ~n14253 & ~n14254;
  assign n14256 = n3457 & n12502;
  assign n14257 = n3542 & n12505;
  assign n14258 = n3606 & n12370;
  assign n14259 = ~n14257 & ~n14258;
  assign n14260 = ~n14256 & n14259;
  assign n14261 = ~n3368 & n14260;
  assign n14262 = n13736 & n14260;
  assign n14263 = ~n14261 & ~n14262;
  assign n14264 =  a[29]  & ~n14263;
  assign n14265 = ~ a[29]  & n14263;
  assign n14266 = ~n14264 & ~n14265;
  assign n14267 = n14255 & ~n14266;
  assign n14268 = ~n14253 & ~n14267;
  assign n14269 = n14062 & n14073;
  assign n14270 = ~n14074 & ~n14269;
  assign n14271 = ~n14268 & n14270;
  assign n14272 = n14268 & ~n14270;
  assign n14273 = ~n14271 & ~n14272;
  assign n14274 = n3884 & n13518;
  assign n14275 = n3967 & n12889;
  assign n14276 = n4046 & n13491;
  assign n14277 = ~n14275 & ~n14276;
  assign n14278 = ~n14274 & n14277;
  assign n14279 = n4050 & n13584;
  assign n14280 = n14278 & ~n14279;
  assign n14281 =  a[26]  & ~n14280;
  assign n14282 =  a[26]  & ~n14281;
  assign n14283 = ~n14280 & ~n14281;
  assign n14284 = ~n14282 & ~n14283;
  assign n14285 = n14273 & ~n14284;
  assign n14286 = ~n14271 & ~n14285;
  assign n14287 = ~n14175 & ~n14286;
  assign n14288 = ~n14172 & ~n14287;
  assign n14289 = ~n14157 & ~n14288;
  assign n14290 = n14157 & n14288;
  assign n14291 = ~n14289 & ~n14290;
  assign n14292 = n4694 & n13633;
  assign n14293 = n4533 & n13597;
  assign n14294 = n4604 & n13630;
  assign n14295 = ~n14293 & ~n14294;
  assign n14296 = ~n14292 & n14295;
  assign n14297 = n4536 & n13929;
  assign n14298 = n14296 & ~n14297;
  assign n14299 =  a[23]  & ~n14298;
  assign n14300 =  a[23]  & ~n14299;
  assign n14301 = ~n14298 & ~n14299;
  assign n14302 = ~n14300 & ~n14301;
  assign n14303 = n14291 & ~n14302;
  assign n14304 = ~n14289 & ~n14303;
  assign n14305 = ~n13438 & ~n13439;
  assign n14306 = n4935 & n13941;
  assign n14307 = ~n14305 & ~n14306;
  assign n14308 = ~n4938 & n14307;
  assign n14309 = n13951 & n14307;
  assign n14310 = ~n14308 & ~n14309;
  assign n14311 =  a[20]  & ~n14310;
  assign n14312 = ~ a[20]  & n14310;
  assign n14313 = ~n14311 & ~n14312;
  assign n14314 = ~n14304 & ~n14313;
  assign n14315 = n14116 & ~n14128;
  assign n14316 = ~n14127 & ~n14128;
  assign n14317 = ~n14315 & ~n14316;
  assign n14318 = n14304 & n14313;
  assign n14319 = ~n14314 & ~n14318;
  assign n14320 = ~n14317 & n14319;
  assign n14321 = ~n14314 & ~n14320;
  assign n14322 = ~n14145 & n14148;
  assign n14323 = ~n14149 & ~n14322;
  assign n14324 = ~n14321 & n14323;
  assign n14325 = ~n14317 & ~n14320;
  assign n14326 = n14319 & ~n14320;
  assign n14327 = ~n14325 & ~n14326;
  assign n14328 = n14291 & ~n14303;
  assign n14329 = ~n14302 & ~n14303;
  assign n14330 = ~n14328 & ~n14329;
  assign n14331 = n14175 & n14286;
  assign n14332 = ~n14287 & ~n14331;
  assign n14333 = n4694 & n13630;
  assign n14334 = n4533 & n13515;
  assign n14335 = n4604 & n13597;
  assign n14336 = ~n14334 & ~n14335;
  assign n14337 = ~n14333 & n14336;
  assign n14338 = n4536 & n13976;
  assign n14339 = n14337 & ~n14338;
  assign n14340 =  a[23]  & ~n14339;
  assign n14341 =  a[23]  & ~n14340;
  assign n14342 = ~n14339 & ~n14340;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = n14332 & ~n14343;
  assign n14345 = n14332 & ~n14344;
  assign n14346 = ~n14343 & ~n14344;
  assign n14347 = ~n14345 & ~n14346;
  assign n14348 = n14273 & ~n14285;
  assign n14349 = ~n14284 & ~n14285;
  assign n14350 = ~n14348 & ~n14349;
  assign n14351 = n14248 & ~n14249;
  assign n14352 = ~n14184 & ~n14249;
  assign n14353 = ~n14351 & ~n14352;
  assign n14354 = n3457 & n12370;
  assign n14355 = n3542 & n12508;
  assign n14356 = n3606 & n12505;
  assign n14357 = ~n14355 & ~n14356;
  assign n14358 = ~n14354 & n14357;
  assign n14359 = n3368 & ~n13748;
  assign n14360 = n14358 & ~n14359;
  assign n14361 =  a[29]  & ~n14360;
  assign n14362 =  a[29]  & ~n14361;
  assign n14363 = ~n14360 & ~n14361;
  assign n14364 = ~n14362 & ~n14363;
  assign n14365 = ~n14353 & ~n14364;
  assign n14366 = ~n14353 & ~n14365;
  assign n14367 = ~n14364 & ~n14365;
  assign n14368 = ~n14366 & ~n14367;
  assign n14369 = ~n14240 & ~n14242;
  assign n14370 = ~n14230 & n14243;
  assign n14371 = ~n14369 & ~n14370;
  assign n14372 = n1271 & n1602;
  assign n14373 = n2698 & n14372;
  assign n14374 = ~n123 & n14373;
  assign n14375 = ~n557 & n14374;
  assign n14376 = ~n571 & n14375;
  assign n14377 = ~n513 & n14376;
  assign n14378 = ~n490 & n14377;
  assign n14379 = ~n302 & n14378;
  assign n14380 = ~n191 & n14379;
  assign n14381 = ~n372 & n14380;
  assign n14382 = ~n278 & n5064;
  assign n14383 = ~n248 & n14382;
  assign n14384 = ~n403 & n14383;
  assign n14385 = ~n164 & n14384;
  assign n14386 = ~n366 & n14385;
  assign n14387 = n1996 & n13114;
  assign n14388 = n4130 & n14387;
  assign n14389 = n2022 & n14388;
  assign n14390 = n14386 & n14389;
  assign n14391 = n2772 & n14390;
  assign n14392 = n6097 & n14391;
  assign n14393 = n14381 & n14392;
  assign n14394 = n2583 & n14393;
  assign n14395 = n1367 & n14394;
  assign n14396 = n1389 & n14395;
  assign n14397 = ~n420 & n14396;
  assign n14398 = ~n281 & n14397;
  assign n14399 = n4294 & n14398;
  assign n14400 = ~n393 & n14399;
  assign n14401 = ~n272 & n14400;
  assign n14402 = ~n672 & n14401;
  assign n14403 = ~n371 & n14402;
  assign n14404 = n1140 & n2210;
  assign n14405 = ~n619 & n14404;
  assign n14406 = ~n157 & n14405;
  assign n14407 = ~n125 & n14406;
  assign n14408 = n889 & n2363;
  assign n14409 = n2544 & n14408;
  assign n14410 = n1085 & n14409;
  assign n14411 = n5746 & n14410;
  assign n14412 = n1119 & n14411;
  assign n14413 = n268 & n14412;
  assign n14414 = n3405 & n14413;
  assign n14415 = n3472 & n14414;
  assign n14416 = n14407 & n14415;
  assign n14417 = n933 & n14416;
  assign n14418 = n4295 & n14417;
  assign n14419 = ~n168 & n14418;
  assign n14420 = ~n400 & n14419;
  assign n14421 = ~n206 & n14420;
  assign n14422 = ~n145 & n14421;
  assign n14423 = ~n14403 & ~n14422;
  assign n14424 = ~n7632 & ~n7983;
  assign n14425 = ~n7291 & n14424;
  assign n14426 = ~n7294 & n14425;
  assign n14427 = ~n13438 & ~n14426;
  assign n14428 =  a[11]  & ~n14427;
  assign n14429 = ~ a[11]  & n14427;
  assign n14430 = ~n14428 & ~n14429;
  assign n14431 = n14403 & n14422;
  assign n14432 = ~n14423 & ~n14431;
  assign n14433 = n14430 & n14432;
  assign n14434 = ~n14423 & ~n14433;
  assign n14435 = n13821 & ~n14434;
  assign n14436 = ~n13821 & n14434;
  assign n14437 = ~n14435 & ~n14436;
  assign n14438 = n3020 & n12516;
  assign n14439 = n3028 & n12519;
  assign n14440 = n3023 & n12522;
  assign n14441 = ~n12655 & ~n12658;
  assign n14442 = ~n12656 & n12659;
  assign n14443 = ~n14441 & ~n14442;
  assign n14444 = n75 & ~n14443;
  assign n14445 = ~n14440 & ~n14444;
  assign n14446 = ~n14439 & n14445;
  assign n14447 = ~n14438 & n14446;
  assign n14448 = n14437 & ~n14447;
  assign n14449 = ~n14435 & ~n14448;
  assign n14450 = ~n14371 & ~n14449;
  assign n14451 = n14371 & n14449;
  assign n14452 = ~n14450 & ~n14451;
  assign n14453 = n12651 & ~n12653;
  assign n14454 = ~n12654 & ~n14453;
  assign n14455 = n75 & n14454;
  assign n14456 = n3020 & n12519;
  assign n14457 = n3023 & n12525;
  assign n14458 = n3028 & n12522;
  assign n14459 = ~n14457 & ~n14458;
  assign n14460 = ~n14456 & n14459;
  assign n14461 = ~n14455 & n14460;
  assign n14462 = ~n14430 & ~n14432;
  assign n14463 = ~n14433 & ~n14462;
  assign n14464 = ~n14461 & n14463;
  assign n14465 = n14463 & ~n14464;
  assign n14466 = ~n14461 & ~n14464;
  assign n14467 = ~n14465 & ~n14466;
  assign n14468 = n1204 & n2154;
  assign n14469 = n665 & n14468;
  assign n14470 = ~n617 & n14469;
  assign n14471 = ~n169 & n14470;
  assign n14472 = ~n667 & n14471;
  assign n14473 = ~n402 & n14472;
  assign n14474 = ~n490 & n14473;
  assign n14475 = ~n374 & n14474;
  assign n14476 = ~n132 & n14475;
  assign n14477 = ~n601 & ~n1101;
  assign n14478 = ~n251 & n14477;
  assign n14479 = ~n270 & n14478;
  assign n14480 = n510 & ~n809;
  assign n14481 = ~n568 & n14480;
  assign n14482 = ~n424 & n14481;
  assign n14483 = n1425 & n3549;
  assign n14484 = n2653 & n14483;
  assign n14485 = n14482 & n14484;
  assign n14486 = n198 & n14485;
  assign n14487 = n1940 & n14486;
  assign n14488 = n14479 & n14487;
  assign n14489 = n1292 & n14488;
  assign n14490 = n1330 & n14489;
  assign n14491 = n827 & n14490;
  assign n14492 = n1380 & n14491;
  assign n14493 = n1269 & n14492;
  assign n14494 = ~n397 & n14493;
  assign n14495 = ~n1246 & n14494;
  assign n14496 = ~n278 & n14495;
  assign n14497 = ~n95 & n14496;
  assign n14498 = ~n125 & n14497;
  assign n14499 = n674 & n1646;
  assign n14500 = n3985 & n14499;
  assign n14501 = n207 & n14500;
  assign n14502 = n14498 & n14501;
  assign n14503 = n4247 & n14502;
  assign n14504 = n14476 & n14503;
  assign n14505 = n622 & n14504;
  assign n14506 = n2739 & n14505;
  assign n14507 = n159 & n14506;
  assign n14508 = n356 & n14507;
  assign n14509 = ~n229 & n14508;
  assign n14510 = ~n620 & n14509;
  assign n14511 = ~n248 & n14510;
  assign n14512 = ~n416 & n14511;
  assign n14513 = ~n237 & n14512;
  assign n14514 = ~n119 & n14513;
  assign n14515 = n14403 & ~n14514;
  assign n14516 = ~n14403 & n14514;
  assign n14517 = ~n118 & n454;
  assign n14518 = ~n165 & n14517;
  assign n14519 = n2348 & n14518;
  assign n14520 = n1576 & n14519;
  assign n14521 = ~n571 & n14520;
  assign n14522 = ~n594 & n14521;
  assign n14523 = ~n132 & n14522;
  assign n14524 = ~n1010 & n14523;
  assign n14525 = ~n270 & n14524;
  assign n14526 = n343 & n13700;
  assign n14527 = n1070 & n14526;
  assign n14528 = n3409 & n14527;
  assign n14529 = ~n1062 & n14528;
  assign n14530 = ~n809 & n14529;
  assign n14531 = ~n331 & n14530;
  assign n14532 = ~n689 & n14531;
  assign n14533 = ~n673 & n14532;
  assign n14534 = ~n474 & n14533;
  assign n14535 = n497 & n1315;
  assign n14536 = n4132 & n14535;
  assign n14537 = n2192 & n14536;
  assign n14538 = n450 & n14537;
  assign n14539 = n227 & n14538;
  assign n14540 = ~n803 & n14539;
  assign n14541 = ~n435 & n14540;
  assign n14542 = ~n461 & n14541;
  assign n14543 = ~n306 & n14542;
  assign n14544 = ~n237 & n14543;
  assign n14545 = n2026 & n2995;
  assign n14546 = n3512 & n14545;
  assign n14547 = n2317 & n14546;
  assign n14548 = n3113 & n14547;
  assign n14549 = n14544 & n14548;
  assign n14550 = n14534 & n14549;
  assign n14551 = n14525 & n14550;
  assign n14552 = n2633 & n14551;
  assign n14553 = n2443 & n14552;
  assign n14554 = n720 & n14553;
  assign n14555 = n356 & n14554;
  assign n14556 = n1180 & n14555;
  assign n14557 = ~n194 & n14556;
  assign n14558 = ~n334 & n14557;
  assign n14559 = ~n125 & n14558;
  assign n14560 = ~n594 & ~n716;
  assign n14561 = ~n331 & n14560;
  assign n14562 = ~n1246 & n14561;
  assign n14563 = ~n289 & n14562;
  assign n14564 = ~n527 & n14563;
  assign n14565 = ~n201 & n14564;
  assign n14566 = n1695 & n2012;
  assign n14567 = n1602 & n14566;
  assign n14568 = n810 & n14567;
  assign n14569 = ~n151 & n14568;
  assign n14570 = ~n286 & n14569;
  assign n14571 = ~n496 & n14570;
  assign n14572 = ~n272 & n14571;
  assign n14573 = n1896 & n2293;
  assign n14574 = n693 & n14573;
  assign n14575 = n5036 & n14574;
  assign n14576 = n1692 & n14575;
  assign n14577 = n13265 & n14576;
  assign n14578 = n14572 & n14577;
  assign n14579 = n1100 & n14578;
  assign n14580 = n120 & n14579;
  assign n14581 = n14565 & n14580;
  assign n14582 = n359 & n14581;
  assign n14583 = ~n427 & n14582;
  assign n14584 = ~n397 & n14583;
  assign n14585 = ~n206 & n14584;
  assign n14586 = ~n505 & n14585;
  assign n14587 = ~n170 & n14586;
  assign n14588 = ~n493 & n14587;
  assign n14589 = ~n14559 & ~n14588;
  assign n14590 = ~n8860 & ~n9331;
  assign n14591 = ~n8418 & n14590;
  assign n14592 = ~n8421 & n14591;
  assign n14593 = ~n13438 & ~n14592;
  assign n14594 =  a[8]  & ~n14593;
  assign n14595 = ~ a[8]  & n14593;
  assign n14596 = ~n14594 & ~n14595;
  assign n14597 = n14559 & n14588;
  assign n14598 = ~n14589 & ~n14597;
  assign n14599 = n14596 & n14598;
  assign n14600 = ~n14589 & ~n14599;
  assign n14601 = n14403 & ~n14600;
  assign n14602 = ~n14403 & n14600;
  assign n14603 = ~n14601 & ~n14602;
  assign n14604 = n3020 & n12525;
  assign n14605 = n3028 & n12528;
  assign n14606 = n3023 & n12531;
  assign n14607 = n12643 & ~n12645;
  assign n14608 = ~n12646 & ~n14607;
  assign n14609 = n75 & n14608;
  assign n14610 = ~n14606 & ~n14609;
  assign n14611 = ~n14605 & n14610;
  assign n14612 = ~n14604 & n14611;
  assign n14613 = n14603 & ~n14612;
  assign n14614 = ~n14601 & ~n14613;
  assign n14615 = ~n14515 & ~n14614;
  assign n14616 = ~n14516 & n14615;
  assign n14617 = ~n14515 & ~n14616;
  assign n14618 = ~n14467 & ~n14617;
  assign n14619 = ~n14464 & ~n14618;
  assign n14620 = ~n14437 & n14447;
  assign n14621 = ~n14448 & ~n14620;
  assign n14622 = ~n14619 & n14621;
  assign n14623 = n14619 & ~n14621;
  assign n14624 = ~n14622 & ~n14623;
  assign n14625 = n3457 & n12508;
  assign n14626 = n3542 & n12511;
  assign n14627 = n3606 & n12513;
  assign n14628 = ~n14626 & ~n14627;
  assign n14629 = ~n14625 & n14628;
  assign n14630 = ~n3368 & n14629;
  assign n14631 = ~n13863 & n14629;
  assign n14632 = ~n14630 & ~n14631;
  assign n14633 =  a[29]  & ~n14632;
  assign n14634 = ~ a[29]  & n14632;
  assign n14635 = ~n14633 & ~n14634;
  assign n14636 = n14624 & ~n14635;
  assign n14637 = ~n14622 & ~n14636;
  assign n14638 = n14452 & ~n14637;
  assign n14639 = ~n14450 & ~n14638;
  assign n14640 = ~n14368 & ~n14639;
  assign n14641 = ~n14365 & ~n14640;
  assign n14642 = ~n14255 & n14266;
  assign n14643 = ~n14267 & ~n14642;
  assign n14644 = ~n14641 & n14643;
  assign n14645 = n14641 & ~n14643;
  assign n14646 = ~n14644 & ~n14645;
  assign n14647 = n3884 & n13491;
  assign n14648 = n3967 & n12769;
  assign n14649 = n4046 & n12889;
  assign n14650 = ~n14648 & ~n14649;
  assign n14651 = ~n14647 & n14650;
  assign n14652 = n4050 & ~n13503;
  assign n14653 = n14651 & ~n14652;
  assign n14654 =  a[26]  & ~n14653;
  assign n14655 =  a[26]  & ~n14654;
  assign n14656 = ~n14653 & ~n14654;
  assign n14657 = ~n14655 & ~n14656;
  assign n14658 = n14646 & ~n14657;
  assign n14659 = ~n14644 & ~n14658;
  assign n14660 = ~n14350 & ~n14659;
  assign n14661 = n14350 & n14659;
  assign n14662 = ~n14660 & ~n14661;
  assign n14663 = n4694 & n13597;
  assign n14664 = n4533 & n13521;
  assign n14665 = n4604 & n13515;
  assign n14666 = ~n14664 & ~n14665;
  assign n14667 = ~n14663 & n14666;
  assign n14668 = n4536 & ~n13612;
  assign n14669 = n14667 & ~n14668;
  assign n14670 =  a[23]  & ~n14669;
  assign n14671 =  a[23]  & ~n14670;
  assign n14672 = ~n14669 & ~n14670;
  assign n14673 = ~n14671 & ~n14672;
  assign n14674 = n14662 & ~n14673;
  assign n14675 = ~n14660 & ~n14674;
  assign n14676 = ~n14347 & ~n14675;
  assign n14677 = ~n14344 & ~n14676;
  assign n14678 = ~n14330 & ~n14677;
  assign n14679 = n14330 & n14677;
  assign n14680 = ~n14678 & ~n14679;
  assign n14681 = n5496 & ~n13438;
  assign n14682 = n4935 & ~n13627;
  assign n14683 = n5407 & n13941;
  assign n14684 = ~n14682 & ~n14683;
  assign n14685 = ~n14681 & n14684;
  assign n14686 = n4938 & n14028;
  assign n14687 = n14685 & ~n14686;
  assign n14688 =  a[20]  & ~n14687;
  assign n14689 =  a[20]  & ~n14688;
  assign n14690 = ~n14687 & ~n14688;
  assign n14691 = ~n14689 & ~n14690;
  assign n14692 = n14680 & ~n14691;
  assign n14693 = ~n14678 & ~n14692;
  assign n14694 = ~n14327 & ~n14693;
  assign n14695 = n14327 & n14693;
  assign n14696 = ~n14694 & ~n14695;
  assign n14697 = n14680 & ~n14692;
  assign n14698 = ~n14691 & ~n14692;
  assign n14699 = ~n14697 & ~n14698;
  assign n14700 = n14662 & ~n14674;
  assign n14701 = ~n14673 & ~n14674;
  assign n14702 = ~n14700 & ~n14701;
  assign n14703 = n14646 & ~n14658;
  assign n14704 = ~n14657 & ~n14658;
  assign n14705 = ~n14703 & ~n14704;
  assign n14706 = n14368 & n14639;
  assign n14707 = ~n14640 & ~n14706;
  assign n14708 = n3884 & n12889;
  assign n14709 = n3967 & n12502;
  assign n14710 = n4046 & n12769;
  assign n14711 = ~n14709 & ~n14710;
  assign n14712 = ~n14708 & n14711;
  assign n14713 = n4050 & n12895;
  assign n14714 = n14712 & ~n14713;
  assign n14715 =  a[26]  & ~n14714;
  assign n14716 =  a[26]  & ~n14715;
  assign n14717 = ~n14714 & ~n14715;
  assign n14718 = ~n14716 & ~n14717;
  assign n14719 = n14707 & ~n14718;
  assign n14720 = n14707 & ~n14719;
  assign n14721 = ~n14718 & ~n14719;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = ~n14452 & n14637;
  assign n14724 = ~n14638 & ~n14723;
  assign n14725 = n3457 & n12505;
  assign n14726 = n3542 & n12513;
  assign n14727 = n3606 & n12508;
  assign n14728 = ~n14726 & ~n14727;
  assign n14729 = ~n14725 & n14728;
  assign n14730 = n3368 & ~n14051;
  assign n14731 = n14729 & ~n14730;
  assign n14732 =  a[29]  & ~n14731;
  assign n14733 =  a[29]  & ~n14732;
  assign n14734 = ~n14731 & ~n14732;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = n14724 & ~n14735;
  assign n14737 = n14724 & ~n14736;
  assign n14738 = ~n14735 & ~n14736;
  assign n14739 = ~n14737 & ~n14738;
  assign n14740 = n3884 & n12769;
  assign n14741 = n3967 & n12370;
  assign n14742 = n4046 & n12502;
  assign n14743 = ~n14741 & ~n14742;
  assign n14744 = ~n14740 & n14743;
  assign n14745 = n4050 & n12999;
  assign n14746 = n14744 & ~n14745;
  assign n14747 =  a[26]  & ~n14746;
  assign n14748 =  a[26]  & ~n14747;
  assign n14749 = ~n14746 & ~n14747;
  assign n14750 = ~n14748 & ~n14749;
  assign n14751 = ~n14739 & ~n14750;
  assign n14752 = ~n14736 & ~n14751;
  assign n14753 = ~n14722 & ~n14752;
  assign n14754 = ~n14719 & ~n14753;
  assign n14755 = ~n14705 & ~n14754;
  assign n14756 = n14705 & n14754;
  assign n14757 = ~n14755 & ~n14756;
  assign n14758 = n4694 & n13515;
  assign n14759 = n4533 & n13518;
  assign n14760 = n4604 & n13521;
  assign n14761 = ~n14759 & ~n14760;
  assign n14762 = ~n14758 & n14761;
  assign n14763 = n4536 & n13541;
  assign n14764 = n14762 & ~n14763;
  assign n14765 =  a[23]  & ~n14764;
  assign n14766 =  a[23]  & ~n14765;
  assign n14767 = ~n14764 & ~n14765;
  assign n14768 = ~n14766 & ~n14767;
  assign n14769 = n14757 & ~n14768;
  assign n14770 = ~n14755 & ~n14769;
  assign n14771 = ~n14702 & ~n14770;
  assign n14772 = n14702 & n14770;
  assign n14773 = ~n14771 & ~n14772;
  assign n14774 = n5496 & ~n13627;
  assign n14775 = n4935 & n13630;
  assign n14776 = n5407 & n13633;
  assign n14777 = ~n14775 & ~n14776;
  assign n14778 = ~n14774 & n14777;
  assign n14779 = n4938 & ~n13654;
  assign n14780 = n14778 & ~n14779;
  assign n14781 =  a[20]  & ~n14780;
  assign n14782 =  a[20]  & ~n14781;
  assign n14783 = ~n14780 & ~n14781;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = n14773 & ~n14784;
  assign n14786 = ~n14771 & ~n14785;
  assign n14787 = n5496 & n13941;
  assign n14788 = n4935 & n13633;
  assign n14789 = n5407 & ~n13627;
  assign n14790 = ~n14788 & ~n14789;
  assign n14791 = ~n14787 & n14790;
  assign n14792 = n4938 & n14136;
  assign n14793 = n14791 & ~n14792;
  assign n14794 =  a[20]  & ~n14793;
  assign n14795 =  a[20]  & ~n14794;
  assign n14796 = ~n14793 & ~n14794;
  assign n14797 = ~n14795 & ~n14796;
  assign n14798 = ~n14786 & ~n14797;
  assign n14799 = n14347 & n14675;
  assign n14800 = ~n14676 & ~n14799;
  assign n14801 = ~n14786 & ~n14798;
  assign n14802 = ~n14797 & ~n14798;
  assign n14803 = ~n14801 & ~n14802;
  assign n14804 = n14800 & ~n14803;
  assign n14805 = ~n14798 & ~n14804;
  assign n14806 = ~n14699 & ~n14805;
  assign n14807 = ~n14699 & ~n14806;
  assign n14808 = ~n14805 & ~n14806;
  assign n14809 = ~n14807 & ~n14808;
  assign n14810 = n14757 & ~n14769;
  assign n14811 = ~n14768 & ~n14769;
  assign n14812 = ~n14810 & ~n14811;
  assign n14813 = n14722 & n14752;
  assign n14814 = ~n14753 & ~n14813;
  assign n14815 = n4694 & n13521;
  assign n14816 = n4533 & n13491;
  assign n14817 = n4604 & n13518;
  assign n14818 = ~n14816 & ~n14817;
  assign n14819 = ~n14815 & n14818;
  assign n14820 = n4536 & ~n13909;
  assign n14821 = n14819 & ~n14820;
  assign n14822 =  a[23]  & ~n14821;
  assign n14823 =  a[23]  & ~n14822;
  assign n14824 = ~n14821 & ~n14822;
  assign n14825 = ~n14823 & ~n14824;
  assign n14826 = n14814 & ~n14825;
  assign n14827 = n14814 & ~n14826;
  assign n14828 = ~n14825 & ~n14826;
  assign n14829 = ~n14827 & ~n14828;
  assign n14830 = ~n14739 & ~n14751;
  assign n14831 = ~n14750 & ~n14751;
  assign n14832 = ~n14830 & ~n14831;
  assign n14833 = ~n14614 & ~n14616;
  assign n14834 = ~n14516 & n14617;
  assign n14835 = ~n14833 & ~n14834;
  assign n14836 = n12647 & ~n12649;
  assign n14837 = ~n12650 & ~n14836;
  assign n14838 = n75 & n14837;
  assign n14839 = n3020 & n12522;
  assign n14840 = n3023 & n12528;
  assign n14841 = n3028 & n12525;
  assign n14842 = ~n14840 & ~n14841;
  assign n14843 = ~n14839 & n14842;
  assign n14844 = ~n14838 & n14843;
  assign n14845 = ~n14835 & ~n14844;
  assign n14846 = ~n14835 & ~n14845;
  assign n14847 = ~n14844 & ~n14845;
  assign n14848 = ~n14846 & ~n14847;
  assign n14849 = n3457 & n12511;
  assign n14850 = n3542 & n12519;
  assign n14851 = n3606 & n12516;
  assign n14852 = ~n14850 & ~n14851;
  assign n14853 = ~n14849 & n14852;
  assign n14854 = ~n3368 & n14853;
  assign n14855 = n14233 & n14853;
  assign n14856 = ~n14854 & ~n14855;
  assign n14857 =  a[29]  & ~n14856;
  assign n14858 = ~ a[29]  & n14856;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = ~n14848 & ~n14859;
  assign n14861 = ~n14845 & ~n14860;
  assign n14862 = ~n14467 & ~n14618;
  assign n14863 = ~n14617 & ~n14618;
  assign n14864 = ~n14862 & ~n14863;
  assign n14865 = ~n14861 & ~n14864;
  assign n14866 = ~n14861 & ~n14865;
  assign n14867 = ~n14864 & ~n14865;
  assign n14868 = ~n14866 & ~n14867;
  assign n14869 = n3457 & n12513;
  assign n14870 = n3542 & n12516;
  assign n14871 = n3606 & n12511;
  assign n14872 = ~n14870 & ~n14871;
  assign n14873 = ~n14869 & n14872;
  assign n14874 = n3368 & n14177;
  assign n14875 = n14873 & ~n14874;
  assign n14876 =  a[29]  & ~n14875;
  assign n14877 =  a[29]  & ~n14876;
  assign n14878 = ~n14875 & ~n14876;
  assign n14879 = ~n14877 & ~n14878;
  assign n14880 = ~n14868 & ~n14879;
  assign n14881 = ~n14865 & ~n14880;
  assign n14882 = ~n14624 & n14635;
  assign n14883 = ~n14636 & ~n14882;
  assign n14884 = ~n14881 & n14883;
  assign n14885 = n14881 & ~n14883;
  assign n14886 = ~n14884 & ~n14885;
  assign n14887 = n3884 & n12502;
  assign n14888 = n3967 & n12505;
  assign n14889 = n4046 & n12370;
  assign n14890 = ~n14888 & ~n14889;
  assign n14891 = ~n14887 & n14890;
  assign n14892 = n4050 & ~n13736;
  assign n14893 = n14891 & ~n14892;
  assign n14894 =  a[26]  & ~n14893;
  assign n14895 =  a[26]  & ~n14894;
  assign n14896 = ~n14893 & ~n14894;
  assign n14897 = ~n14895 & ~n14896;
  assign n14898 = n14886 & ~n14897;
  assign n14899 = ~n14884 & ~n14898;
  assign n14900 = ~n14832 & ~n14899;
  assign n14901 = n14832 & n14899;
  assign n14902 = ~n14900 & ~n14901;
  assign n14903 = n4694 & n13518;
  assign n14904 = n4533 & n12889;
  assign n14905 = n4604 & n13491;
  assign n14906 = ~n14904 & ~n14905;
  assign n14907 = ~n14903 & n14906;
  assign n14908 = n4536 & n13584;
  assign n14909 = n14907 & ~n14908;
  assign n14910 =  a[23]  & ~n14909;
  assign n14911 =  a[23]  & ~n14910;
  assign n14912 = ~n14909 & ~n14910;
  assign n14913 = ~n14911 & ~n14912;
  assign n14914 = n14902 & ~n14913;
  assign n14915 = ~n14900 & ~n14914;
  assign n14916 = ~n14829 & ~n14915;
  assign n14917 = ~n14826 & ~n14916;
  assign n14918 = ~n14812 & ~n14917;
  assign n14919 = n14812 & n14917;
  assign n14920 = ~n14918 & ~n14919;
  assign n14921 = n5496 & n13633;
  assign n14922 = n4935 & n13597;
  assign n14923 = n5407 & n13630;
  assign n14924 = ~n14922 & ~n14923;
  assign n14925 = ~n14921 & n14924;
  assign n14926 = n4938 & n13929;
  assign n14927 = n14925 & ~n14926;
  assign n14928 =  a[20]  & ~n14927;
  assign n14929 =  a[20]  & ~n14928;
  assign n14930 = ~n14927 & ~n14928;
  assign n14931 = ~n14929 & ~n14930;
  assign n14932 = n14920 & ~n14931;
  assign n14933 = ~n14918 & ~n14932;
  assign n14934 = ~n13438 & ~n13717;
  assign n14935 = n5663 & n13941;
  assign n14936 = ~n14934 & ~n14935;
  assign n14937 = ~n5666 & n14936;
  assign n14938 = n13951 & n14936;
  assign n14939 = ~n14937 & ~n14938;
  assign n14940 =  a[17]  & ~n14939;
  assign n14941 = ~ a[17]  & n14939;
  assign n14942 = ~n14940 & ~n14941;
  assign n14943 = ~n14933 & ~n14942;
  assign n14944 = n14773 & ~n14785;
  assign n14945 = ~n14784 & ~n14785;
  assign n14946 = ~n14944 & ~n14945;
  assign n14947 = n14933 & n14942;
  assign n14948 = ~n14943 & ~n14947;
  assign n14949 = ~n14946 & n14948;
  assign n14950 = ~n14943 & ~n14949;
  assign n14951 = ~n14800 & n14803;
  assign n14952 = ~n14804 & ~n14951;
  assign n14953 = ~n14950 & n14952;
  assign n14954 = ~n14946 & ~n14949;
  assign n14955 = n14948 & ~n14949;
  assign n14956 = ~n14954 & ~n14955;
  assign n14957 = n14920 & ~n14932;
  assign n14958 = ~n14931 & ~n14932;
  assign n14959 = ~n14957 & ~n14958;
  assign n14960 = n14829 & n14915;
  assign n14961 = ~n14916 & ~n14960;
  assign n14962 = n5496 & n13630;
  assign n14963 = n4935 & n13515;
  assign n14964 = n5407 & n13597;
  assign n14965 = ~n14963 & ~n14964;
  assign n14966 = ~n14962 & n14965;
  assign n14967 = n4938 & n13976;
  assign n14968 = n14966 & ~n14967;
  assign n14969 =  a[20]  & ~n14968;
  assign n14970 =  a[20]  & ~n14969;
  assign n14971 = ~n14968 & ~n14969;
  assign n14972 = ~n14970 & ~n14971;
  assign n14973 = n14961 & ~n14972;
  assign n14974 = n14961 & ~n14973;
  assign n14975 = ~n14972 & ~n14973;
  assign n14976 = ~n14974 & ~n14975;
  assign n14977 = n14902 & ~n14914;
  assign n14978 = ~n14913 & ~n14914;
  assign n14979 = ~n14977 & ~n14978;
  assign n14980 = n14886 & ~n14898;
  assign n14981 = ~n14897 & ~n14898;
  assign n14982 = ~n14980 & ~n14981;
  assign n14983 = ~n14868 & ~n14880;
  assign n14984 = ~n14879 & ~n14880;
  assign n14985 = ~n14983 & ~n14984;
  assign n14986 = n3884 & n12370;
  assign n14987 = n3967 & n12508;
  assign n14988 = n4046 & n12505;
  assign n14989 = ~n14987 & ~n14988;
  assign n14990 = ~n14986 & n14989;
  assign n14991 = n4050 & ~n13748;
  assign n14992 = n14990 & ~n14991;
  assign n14993 =  a[26]  & ~n14992;
  assign n14994 =  a[26]  & ~n14993;
  assign n14995 = ~n14992 & ~n14993;
  assign n14996 = ~n14994 & ~n14995;
  assign n14997 = ~n14985 & ~n14996;
  assign n14998 = ~n14985 & ~n14997;
  assign n14999 = ~n14996 & ~n14997;
  assign n15000 = ~n14998 & ~n14999;
  assign n15001 = ~n12639 & ~n12642;
  assign n15002 = ~n12640 & n12643;
  assign n15003 = ~n15001 & ~n15002;
  assign n15004 = n75 & ~n15003;
  assign n15005 = n3020 & n12528;
  assign n15006 = n3023 & n12534;
  assign n15007 = n3028 & n12531;
  assign n15008 = ~n15006 & ~n15007;
  assign n15009 = ~n15005 & n15008;
  assign n15010 = ~n15004 & n15009;
  assign n15011 = ~n667 & n1139;
  assign n15012 = ~n886 & n15011;
  assign n15013 = n256 & n5173;
  assign n15014 = n15012 & n15013;
  assign n15015 = n2093 & n15014;
  assign n15016 = n1958 & n15015;
  assign n15017 = n3565 & n15016;
  assign n15018 = n2738 & n15017;
  assign n15019 = n187 & n15018;
  assign n15020 = n2170 & n15019;
  assign n15021 = n471 & n15020;
  assign n15022 = n1857 & n15021;
  assign n15023 = ~n427 & n15022;
  assign n15024 = ~n289 & n15023;
  assign n15025 = ~n281 & n15024;
  assign n15026 = ~n557 & n15025;
  assign n15027 = ~n237 & n15026;
  assign n15028 = ~n201 & n15027;
  assign n15029 = n14559 & ~n15028;
  assign n15030 = ~n14559 & n15028;
  assign n15031 = n11053 & n11054;
  assign n15032 = ~n13438 & ~n15031;
  assign n15033 =  a[2]  & ~n15032;
  assign n15034 = ~ a[2]  & n15032;
  assign n15035 = ~n15033 & ~n15034;
  assign n15036 = n1738 & n3645;
  assign n15037 = n1070 & n15036;
  assign n15038 = n3548 & n15037;
  assign n15039 = n439 & n15038;
  assign n15040 = n508 & n15039;
  assign n15041 = ~n168 & n15040;
  assign n15042 = ~n402 & n15041;
  assign n15043 = ~n961 & n15042;
  assign n15044 = ~n170 & n15043;
  assign n15045 = ~n1010 & n15044;
  assign n15046 = ~n489 & n15045;
  assign n15047 = ~n771 & n15046;
  assign n15048 = n2651 & n14479;
  assign n15049 = ~n301 & n15048;
  assign n15050 = ~n229 & n15049;
  assign n15051 = n3194 & n13827;
  assign n15052 = n370 & n15051;
  assign n15053 = n2241 & n15052;
  assign n15054 = n15050 & n15053;
  assign n15055 = n12810 & n15054;
  assign n15056 = n2591 & n15055;
  assign n15057 = n294 & n15056;
  assign n15058 = n1781 & n15057;
  assign n15059 = n15047 & n15058;
  assign n15060 = n1389 & n15059;
  assign n15061 = ~n417 & n15060;
  assign n15062 = n137 & n3192;
  assign n15063 = n6102 & n15062;
  assign n15064 = n6667 & n15063;
  assign n15065 = n14381 & n15064;
  assign n15066 = n12404 & n15065;
  assign n15067 = n15061 & n15066;
  assign n15068 = n1523 & n15067;
  assign n15069 = n247 & n15068;
  assign n15070 = n3252 & n15069;
  assign n15071 = ~n620 & n15070;
  assign n15072 = ~n352 & n15071;
  assign n15073 = ~n118 & n15072;
  assign n15074 = ~n532 & n15073;
  assign n15075 = n15035 & ~n15074;
  assign n15076 = ~n71 & ~n10434;
  assign n15077 = ~n9867 & n15076;
  assign n15078 = ~n9870 & n15077;
  assign n15079 = ~n13438 & ~n15078;
  assign n15080 = ~ a[5]  & n15079;
  assign n15081 = n15035 & n15074;
  assign n15082 = ~n15035 & ~n15074;
  assign n15083 = ~n15081 & ~n15082;
  assign n15084 =  a[5]  & ~n15079;
  assign n15085 = ~n15083 & ~n15084;
  assign n15086 = ~n15080 & n15085;
  assign n15087 = ~n15075 & ~n15086;
  assign n15088 = n14559 & ~n15087;
  assign n15089 = ~n14559 & n15087;
  assign n15090 = ~n15088 & ~n15089;
  assign n15091 = n3020 & n12534;
  assign n15092 = n3028 & n12537;
  assign n15093 = n3023 & n12540;
  assign n15094 = ~n12631 & ~n12634;
  assign n15095 = ~n12632 & n12635;
  assign n15096 = ~n15094 & ~n15095;
  assign n15097 = n75 & ~n15096;
  assign n15098 = ~n15093 & ~n15097;
  assign n15099 = ~n15092 & n15098;
  assign n15100 = ~n15091 & n15099;
  assign n15101 = n15090 & ~n15100;
  assign n15102 = ~n15088 & ~n15101;
  assign n15103 = ~n15029 & ~n15102;
  assign n15104 = ~n15030 & n15103;
  assign n15105 = ~n15029 & ~n15104;
  assign n15106 = ~n14596 & ~n14598;
  assign n15107 = ~n14599 & ~n15106;
  assign n15108 = ~n15105 & n15107;
  assign n15109 = n15105 & ~n15107;
  assign n15110 = ~n15108 & ~n15109;
  assign n15111 = ~n15010 & n15110;
  assign n15112 = ~n15108 & ~n15111;
  assign n15113 = ~n14603 & n14612;
  assign n15114 = ~n14613 & ~n15113;
  assign n15115 = ~n15112 & n15114;
  assign n15116 = n15112 & ~n15114;
  assign n15117 = ~n15115 & ~n15116;
  assign n15118 = n3457 & n12516;
  assign n15119 = n3542 & n12522;
  assign n15120 = n3606 & n12519;
  assign n15121 = ~n15119 & ~n15120;
  assign n15122 = ~n15118 & n15121;
  assign n15123 = ~n3368 & n15122;
  assign n15124 = n14443 & n15122;
  assign n15125 = ~n15123 & ~n15124;
  assign n15126 =  a[29]  & ~n15125;
  assign n15127 = ~ a[29]  & n15125;
  assign n15128 = ~n15126 & ~n15127;
  assign n15129 = n15117 & ~n15128;
  assign n15130 = ~n15115 & ~n15129;
  assign n15131 = n14848 & n14859;
  assign n15132 = ~n14860 & ~n15131;
  assign n15133 = ~n15130 & n15132;
  assign n15134 = n15130 & ~n15132;
  assign n15135 = ~n15133 & ~n15134;
  assign n15136 = n3884 & n12505;
  assign n15137 = n3967 & n12513;
  assign n15138 = n4046 & n12508;
  assign n15139 = ~n15137 & ~n15138;
  assign n15140 = ~n15136 & n15139;
  assign n15141 = n4050 & ~n14051;
  assign n15142 = n15140 & ~n15141;
  assign n15143 =  a[26]  & ~n15142;
  assign n15144 =  a[26]  & ~n15143;
  assign n15145 = ~n15142 & ~n15143;
  assign n15146 = ~n15144 & ~n15145;
  assign n15147 = n15135 & ~n15146;
  assign n15148 = ~n15133 & ~n15147;
  assign n15149 = ~n15000 & ~n15148;
  assign n15150 = ~n14997 & ~n15149;
  assign n15151 = ~n14982 & ~n15150;
  assign n15152 = n14982 & n15150;
  assign n15153 = ~n15151 & ~n15152;
  assign n15154 = n4694 & n13491;
  assign n15155 = n4533 & n12769;
  assign n15156 = n4604 & n12889;
  assign n15157 = ~n15155 & ~n15156;
  assign n15158 = ~n15154 & n15157;
  assign n15159 = n4536 & ~n13503;
  assign n15160 = n15158 & ~n15159;
  assign n15161 =  a[23]  & ~n15160;
  assign n15162 =  a[23]  & ~n15161;
  assign n15163 = ~n15160 & ~n15161;
  assign n15164 = ~n15162 & ~n15163;
  assign n15165 = n15153 & ~n15164;
  assign n15166 = ~n15151 & ~n15165;
  assign n15167 = ~n14979 & ~n15166;
  assign n15168 = n14979 & n15166;
  assign n15169 = ~n15167 & ~n15168;
  assign n15170 = n5496 & n13597;
  assign n15171 = n4935 & n13521;
  assign n15172 = n5407 & n13515;
  assign n15173 = ~n15171 & ~n15172;
  assign n15174 = ~n15170 & n15173;
  assign n15175 = n4938 & ~n13612;
  assign n15176 = n15174 & ~n15175;
  assign n15177 =  a[20]  & ~n15176;
  assign n15178 =  a[20]  & ~n15177;
  assign n15179 = ~n15176 & ~n15177;
  assign n15180 = ~n15178 & ~n15179;
  assign n15181 = n15169 & ~n15180;
  assign n15182 = ~n15167 & ~n15181;
  assign n15183 = ~n14976 & ~n15182;
  assign n15184 = ~n14973 & ~n15183;
  assign n15185 = ~n14959 & ~n15184;
  assign n15186 = n14959 & n15184;
  assign n15187 = ~n15185 & ~n15186;
  assign n15188 = n6233 & ~n13438;
  assign n15189 = n5663 & ~n13627;
  assign n15190 = n5939 & n13941;
  assign n15191 = ~n15189 & ~n15190;
  assign n15192 = ~n15188 & n15191;
  assign n15193 = n5666 & n14028;
  assign n15194 = n15192 & ~n15193;
  assign n15195 =  a[17]  & ~n15194;
  assign n15196 =  a[17]  & ~n15195;
  assign n15197 = ~n15194 & ~n15195;
  assign n15198 = ~n15196 & ~n15197;
  assign n15199 = n15187 & ~n15198;
  assign n15200 = ~n15185 & ~n15199;
  assign n15201 = ~n14956 & ~n15200;
  assign n15202 = n14956 & n15200;
  assign n15203 = ~n15201 & ~n15202;
  assign n15204 = n15187 & ~n15199;
  assign n15205 = ~n15198 & ~n15199;
  assign n15206 = ~n15204 & ~n15205;
  assign n15207 = n15169 & ~n15181;
  assign n15208 = ~n15180 & ~n15181;
  assign n15209 = ~n15207 & ~n15208;
  assign n15210 = n15153 & ~n15165;
  assign n15211 = ~n15164 & ~n15165;
  assign n15212 = ~n15210 & ~n15211;
  assign n15213 = n15000 & n15148;
  assign n15214 = ~n15149 & ~n15213;
  assign n15215 = n4694 & n12889;
  assign n15216 = n4533 & n12502;
  assign n15217 = n4604 & n12769;
  assign n15218 = ~n15216 & ~n15217;
  assign n15219 = ~n15215 & n15218;
  assign n15220 = n4536 & n12895;
  assign n15221 = n15219 & ~n15220;
  assign n15222 =  a[23]  & ~n15221;
  assign n15223 =  a[23]  & ~n15222;
  assign n15224 = ~n15221 & ~n15222;
  assign n15225 = ~n15223 & ~n15224;
  assign n15226 = n15214 & ~n15225;
  assign n15227 = n15214 & ~n15226;
  assign n15228 = ~n15225 & ~n15226;
  assign n15229 = ~n15227 & ~n15228;
  assign n15230 = n15135 & ~n15147;
  assign n15231 = ~n15146 & ~n15147;
  assign n15232 = ~n15230 & ~n15231;
  assign n15233 = n15110 & ~n15111;
  assign n15234 = ~n15010 & ~n15111;
  assign n15235 = ~n15233 & ~n15234;
  assign n15236 = n3457 & n12519;
  assign n15237 = n3542 & n12525;
  assign n15238 = n3606 & n12522;
  assign n15239 = ~n15237 & ~n15238;
  assign n15240 = ~n15236 & n15239;
  assign n15241 = n3368 & n14454;
  assign n15242 = n15240 & ~n15241;
  assign n15243 =  a[29]  & ~n15242;
  assign n15244 =  a[29]  & ~n15243;
  assign n15245 = ~n15242 & ~n15243;
  assign n15246 = ~n15244 & ~n15245;
  assign n15247 = ~n15235 & ~n15246;
  assign n15248 = ~n15235 & ~n15247;
  assign n15249 = ~n15246 & ~n15247;
  assign n15250 = ~n15248 & ~n15249;
  assign n15251 = ~n15102 & ~n15104;
  assign n15252 = ~n15030 & n15105;
  assign n15253 = ~n15251 & ~n15252;
  assign n15254 = n12635 & ~n12637;
  assign n15255 = ~n12638 & ~n15254;
  assign n15256 = n75 & n15255;
  assign n15257 = n3020 & n12531;
  assign n15258 = n3023 & n12537;
  assign n15259 = n3028 & n12534;
  assign n15260 = ~n15258 & ~n15259;
  assign n15261 = ~n15257 & n15260;
  assign n15262 = ~n15256 & n15261;
  assign n15263 = ~n15253 & ~n15262;
  assign n15264 = ~n15253 & ~n15263;
  assign n15265 = ~n15262 & ~n15263;
  assign n15266 = ~n15264 & ~n15265;
  assign n15267 = n1185 & n2349;
  assign n15268 = n1894 & n15267;
  assign n15269 = n3743 & n15268;
  assign n15270 = n3675 & n15269;
  assign n15271 = n5785 & n15270;
  assign n15272 = n2778 & n15271;
  assign n15273 = n1180 & n15272;
  assign n15274 = ~n469 & n15273;
  assign n15275 = ~n1101 & n15274;
  assign n15276 = ~n513 & n15275;
  assign n15277 = ~n298 & n15276;
  assign n15278 = ~n372 & n15277;
  assign n15279 = ~n157 & n15278;
  assign n15280 = ~n1104 & n15279;
  assign n15281 = ~n592 & n15280;
  assign n15282 = ~n295 & n15281;
  assign n15283 = ~n525 & n15282;
  assign n15284 = ~n15035 & ~n15283;
  assign n15285 = n634 & n13774;
  assign n15286 = ~n328 & n15285;
  assign n15287 = n13012 & n15286;
  assign n15288 = n1709 & n15287;
  assign n15289 = n15061 & n15288;
  assign n15290 = n503 & n15289;
  assign n15291 = n512 & n15290;
  assign n15292 = n1915 & n15291;
  assign n15293 = n1183 & n15292;
  assign n15294 = n285 & n15293;
  assign n15295 = n730 & n15294;
  assign n15296 = n1783 & n15295;
  assign n15297 = n202 & n15296;
  assign n15298 = n4101 & n15297;
  assign n15299 = ~n746 & n15298;
  assign n15300 = ~n239 & n15299;
  assign n15301 = ~n192 & n15300;
  assign n15302 = ~n453 & n15301;
  assign n15303 = ~n883 & n15302;
  assign n15304 = ~n886 & n15303;
  assign n15305 = ~n337 & n15304;
  assign n15306 = ~n15035 & ~n15305;
  assign n15307 = n1557 & n2209;
  assign n15308 = ~n420 & n15307;
  assign n15309 = ~n278 & n15308;
  assign n15310 = ~n435 & n15309;
  assign n15311 = ~n589 & n15310;
  assign n15312 = ~n569 & n15311;
  assign n15313 = n365 & n1329;
  assign n15314 = n2468 & n15313;
  assign n15315 = n12431 & n15314;
  assign n15316 = n5085 & n15315;
  assign n15317 = n1725 & n15316;
  assign n15318 = n15312 & n15317;
  assign n15319 = n2346 & n15318;
  assign n15320 = ~n151 & n15319;
  assign n15321 = ~n275 & n15320;
  assign n15322 = ~n438 & n15321;
  assign n15323 = ~n1203 & n15322;
  assign n15324 = ~n623 & n15323;
  assign n15325 = n1692 & n15324;
  assign n15326 = ~n354 & n15325;
  assign n15327 = ~n168 & n15326;
  assign n15328 = ~n296 & n15327;
  assign n15329 = ~n1104 & n15328;
  assign n15330 = ~n532 & n15329;
  assign n15331 = ~n1306 & n3380;
  assign n15332 = ~n746 & n15331;
  assign n15333 = ~n232 & n15332;
  assign n15334 = ~n152 & n15333;
  assign n15335 = ~n203 & n15334;
  assign n15336 = ~n245 & n15335;
  assign n15337 = ~n932 & n15336;
  assign n15338 = n475 & n1530;
  assign n15339 = n2809 & n15338;
  assign n15340 = n1759 & n15339;
  assign n15341 = n15337 & n15340;
  assign n15342 = n12973 & n15341;
  assign n15343 = n15330 & n15342;
  assign n15344 = n14479 & n15343;
  assign n15345 = n1237 & n15344;
  assign n15346 = ~n111 & n15345;
  assign n15347 = ~n150 & n15346;
  assign n15348 = ~n571 & n15347;
  assign n15349 = ~n118 & n15348;
  assign n15350 = ~n107 & n15349;
  assign n15351 = ~n286 & n15350;
  assign n15352 = ~n592 & n15351;
  assign n15353 = ~n15035 & ~n15352;
  assign n15354 = ~n12615 & ~n12618;
  assign n15355 = ~n12616 & n12619;
  assign n15356 = ~n15354 & ~n15355;
  assign n15357 = n75 & ~n15356;
  assign n15358 = n3020 & n12546;
  assign n15359 = n3023 & n12552;
  assign n15360 = n3028 & n12549;
  assign n15361 = ~n15359 & ~n15360;
  assign n15362 = ~n15358 & n15361;
  assign n15363 = ~n15357 & n15362;
  assign n15364 = n15035 & n15352;
  assign n15365 = ~n15363 & ~n15364;
  assign n15366 = ~n15353 & n15365;
  assign n15367 = ~n15353 & ~n15366;
  assign n15368 = n15035 & n15305;
  assign n15369 = ~n15367 & ~n15368;
  assign n15370 = ~n15306 & n15369;
  assign n15371 = ~n15306 & ~n15370;
  assign n15372 = n15035 & n15283;
  assign n15373 = ~n15371 & ~n15372;
  assign n15374 = ~n15284 & n15373;
  assign n15375 = ~n15284 & ~n15374;
  assign n15376 = ~n15083 & ~n15086;
  assign n15377 = ~n15084 & ~n15086;
  assign n15378 = ~n15080 & n15377;
  assign n15379 = ~n15376 & ~n15378;
  assign n15380 = ~n15375 & n15379;
  assign n15381 = n15375 & ~n15379;
  assign n15382 = ~n15380 & ~n15381;
  assign n15383 = ~n12627 & ~n12630;
  assign n15384 = ~n12628 & n12631;
  assign n15385 = ~n15383 & ~n15384;
  assign n15386 = n75 & ~n15385;
  assign n15387 = n3020 & n12537;
  assign n15388 = n3023 & n12543;
  assign n15389 = n3028 & n12540;
  assign n15390 = ~n15388 & ~n15389;
  assign n15391 = ~n15387 & n15390;
  assign n15392 = ~n15386 & n15391;
  assign n15393 = ~n15382 & ~n15392;
  assign n15394 = ~n15375 & ~n15379;
  assign n15395 = ~n15393 & ~n15394;
  assign n15396 = ~n15090 & n15100;
  assign n15397 = ~n15101 & ~n15396;
  assign n15398 = ~n15395 & n15397;
  assign n15399 = n15395 & ~n15397;
  assign n15400 = ~n15398 & ~n15399;
  assign n15401 = n3457 & n12525;
  assign n15402 = n3542 & n12531;
  assign n15403 = n3606 & n12528;
  assign n15404 = ~n15402 & ~n15403;
  assign n15405 = ~n15401 & n15404;
  assign n15406 = ~n3368 & n15405;
  assign n15407 = ~n14608 & n15405;
  assign n15408 = ~n15406 & ~n15407;
  assign n15409 =  a[29]  & ~n15408;
  assign n15410 = ~ a[29]  & n15408;
  assign n15411 = ~n15409 & ~n15410;
  assign n15412 = n15400 & ~n15411;
  assign n15413 = ~n15398 & ~n15412;
  assign n15414 = ~n15266 & ~n15413;
  assign n15415 = ~n15263 & ~n15414;
  assign n15416 = ~n15250 & ~n15415;
  assign n15417 = ~n15247 & ~n15416;
  assign n15418 = ~n15117 & n15128;
  assign n15419 = ~n15129 & ~n15418;
  assign n15420 = ~n15417 & n15419;
  assign n15421 = n15417 & ~n15419;
  assign n15422 = ~n15420 & ~n15421;
  assign n15423 = n3884 & n12508;
  assign n15424 = n3967 & n12511;
  assign n15425 = n4046 & n12513;
  assign n15426 = ~n15424 & ~n15425;
  assign n15427 = ~n15423 & n15426;
  assign n15428 = n4050 & n13863;
  assign n15429 = n15427 & ~n15428;
  assign n15430 =  a[26]  & ~n15429;
  assign n15431 =  a[26]  & ~n15430;
  assign n15432 = ~n15429 & ~n15430;
  assign n15433 = ~n15431 & ~n15432;
  assign n15434 = n15422 & ~n15433;
  assign n15435 = ~n15420 & ~n15434;
  assign n15436 = ~n15232 & ~n15435;
  assign n15437 = n15232 & n15435;
  assign n15438 = ~n15436 & ~n15437;
  assign n15439 = n4694 & n12769;
  assign n15440 = n4533 & n12370;
  assign n15441 = n4604 & n12502;
  assign n15442 = ~n15440 & ~n15441;
  assign n15443 = ~n15439 & n15442;
  assign n15444 = n4536 & n12999;
  assign n15445 = n15443 & ~n15444;
  assign n15446 =  a[23]  & ~n15445;
  assign n15447 =  a[23]  & ~n15446;
  assign n15448 = ~n15445 & ~n15446;
  assign n15449 = ~n15447 & ~n15448;
  assign n15450 = n15438 & ~n15449;
  assign n15451 = ~n15436 & ~n15450;
  assign n15452 = ~n15229 & ~n15451;
  assign n15453 = ~n15226 & ~n15452;
  assign n15454 = ~n15212 & ~n15453;
  assign n15455 = n15212 & n15453;
  assign n15456 = ~n15454 & ~n15455;
  assign n15457 = n5496 & n13515;
  assign n15458 = n4935 & n13518;
  assign n15459 = n5407 & n13521;
  assign n15460 = ~n15458 & ~n15459;
  assign n15461 = ~n15457 & n15460;
  assign n15462 = n4938 & n13541;
  assign n15463 = n15461 & ~n15462;
  assign n15464 =  a[20]  & ~n15463;
  assign n15465 =  a[20]  & ~n15464;
  assign n15466 = ~n15463 & ~n15464;
  assign n15467 = ~n15465 & ~n15466;
  assign n15468 = n15456 & ~n15467;
  assign n15469 = ~n15454 & ~n15468;
  assign n15470 = ~n15209 & ~n15469;
  assign n15471 = n15209 & n15469;
  assign n15472 = ~n15470 & ~n15471;
  assign n15473 = n6233 & ~n13627;
  assign n15474 = n5663 & n13630;
  assign n15475 = n5939 & n13633;
  assign n15476 = ~n15474 & ~n15475;
  assign n15477 = ~n15473 & n15476;
  assign n15478 = n5666 & ~n13654;
  assign n15479 = n15477 & ~n15478;
  assign n15480 =  a[17]  & ~n15479;
  assign n15481 =  a[17]  & ~n15480;
  assign n15482 = ~n15479 & ~n15480;
  assign n15483 = ~n15481 & ~n15482;
  assign n15484 = n15472 & ~n15483;
  assign n15485 = ~n15470 & ~n15484;
  assign n15486 = n6233 & n13941;
  assign n15487 = n5663 & n13633;
  assign n15488 = n5939 & ~n13627;
  assign n15489 = ~n15487 & ~n15488;
  assign n15490 = ~n15486 & n15489;
  assign n15491 = n5666 & n14136;
  assign n15492 = n15490 & ~n15491;
  assign n15493 =  a[17]  & ~n15492;
  assign n15494 =  a[17]  & ~n15493;
  assign n15495 = ~n15492 & ~n15493;
  assign n15496 = ~n15494 & ~n15495;
  assign n15497 = ~n15485 & ~n15496;
  assign n15498 = n14976 & n15182;
  assign n15499 = ~n15183 & ~n15498;
  assign n15500 = ~n15485 & ~n15497;
  assign n15501 = ~n15496 & ~n15497;
  assign n15502 = ~n15500 & ~n15501;
  assign n15503 = n15499 & ~n15502;
  assign n15504 = ~n15497 & ~n15503;
  assign n15505 = ~n15206 & ~n15504;
  assign n15506 = ~n15206 & ~n15505;
  assign n15507 = ~n15504 & ~n15505;
  assign n15508 = ~n15506 & ~n15507;
  assign n15509 = n15456 & ~n15468;
  assign n15510 = ~n15467 & ~n15468;
  assign n15511 = ~n15509 & ~n15510;
  assign n15512 = n15229 & n15451;
  assign n15513 = ~n15452 & ~n15512;
  assign n15514 = n5496 & n13521;
  assign n15515 = n4935 & n13491;
  assign n15516 = n5407 & n13518;
  assign n15517 = ~n15515 & ~n15516;
  assign n15518 = ~n15514 & n15517;
  assign n15519 = n4938 & ~n13909;
  assign n15520 = n15518 & ~n15519;
  assign n15521 =  a[20]  & ~n15520;
  assign n15522 =  a[20]  & ~n15521;
  assign n15523 = ~n15520 & ~n15521;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = n15513 & ~n15524;
  assign n15526 = n15513 & ~n15525;
  assign n15527 = ~n15524 & ~n15525;
  assign n15528 = ~n15526 & ~n15527;
  assign n15529 = n15438 & ~n15450;
  assign n15530 = ~n15449 & ~n15450;
  assign n15531 = ~n15529 & ~n15530;
  assign n15532 = n15422 & ~n15434;
  assign n15533 = ~n15433 & ~n15434;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = n15250 & n15415;
  assign n15536 = ~n15416 & ~n15535;
  assign n15537 = n3884 & n12513;
  assign n15538 = n3967 & n12516;
  assign n15539 = n4046 & n12511;
  assign n15540 = ~n15538 & ~n15539;
  assign n15541 = ~n15537 & n15540;
  assign n15542 = n4050 & n14177;
  assign n15543 = n15541 & ~n15542;
  assign n15544 =  a[26]  & ~n15543;
  assign n15545 =  a[26]  & ~n15544;
  assign n15546 = ~n15543 & ~n15544;
  assign n15547 = ~n15545 & ~n15546;
  assign n15548 = n15536 & ~n15547;
  assign n15549 = n15536 & ~n15548;
  assign n15550 = ~n15547 & ~n15548;
  assign n15551 = ~n15549 & ~n15550;
  assign n15552 = n15266 & n15413;
  assign n15553 = ~n15414 & ~n15552;
  assign n15554 = n3457 & n12522;
  assign n15555 = n3542 & n12528;
  assign n15556 = n3606 & n12525;
  assign n15557 = ~n15555 & ~n15556;
  assign n15558 = ~n15554 & n15557;
  assign n15559 = n3368 & n14837;
  assign n15560 = n15558 & ~n15559;
  assign n15561 =  a[29]  & ~n15560;
  assign n15562 =  a[29]  & ~n15561;
  assign n15563 = ~n15560 & ~n15561;
  assign n15564 = ~n15562 & ~n15563;
  assign n15565 = n15553 & ~n15564;
  assign n15566 = n15553 & ~n15565;
  assign n15567 = ~n15564 & ~n15565;
  assign n15568 = ~n15566 & ~n15567;
  assign n15569 = n3884 & n12511;
  assign n15570 = n3967 & n12519;
  assign n15571 = n4046 & n12516;
  assign n15572 = ~n15570 & ~n15571;
  assign n15573 = ~n15569 & n15572;
  assign n15574 = n4050 & ~n14233;
  assign n15575 = n15573 & ~n15574;
  assign n15576 =  a[26]  & ~n15575;
  assign n15577 =  a[26]  & ~n15576;
  assign n15578 = ~n15575 & ~n15576;
  assign n15579 = ~n15577 & ~n15578;
  assign n15580 = ~n15568 & ~n15579;
  assign n15581 = ~n15565 & ~n15580;
  assign n15582 = ~n15551 & ~n15581;
  assign n15583 = ~n15548 & ~n15582;
  assign n15584 = ~n15534 & ~n15583;
  assign n15585 = n15534 & n15583;
  assign n15586 = ~n15584 & ~n15585;
  assign n15587 = n4694 & n12502;
  assign n15588 = n4533 & n12505;
  assign n15589 = n4604 & n12370;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = ~n15587 & n15590;
  assign n15592 = n4536 & ~n13736;
  assign n15593 = n15591 & ~n15592;
  assign n15594 =  a[23]  & ~n15593;
  assign n15595 =  a[23]  & ~n15594;
  assign n15596 = ~n15593 & ~n15594;
  assign n15597 = ~n15595 & ~n15596;
  assign n15598 = n15586 & ~n15597;
  assign n15599 = ~n15584 & ~n15598;
  assign n15600 = ~n15531 & ~n15599;
  assign n15601 = n15531 & n15599;
  assign n15602 = ~n15600 & ~n15601;
  assign n15603 = n5496 & n13518;
  assign n15604 = n4935 & n12889;
  assign n15605 = n5407 & n13491;
  assign n15606 = ~n15604 & ~n15605;
  assign n15607 = ~n15603 & n15606;
  assign n15608 = n4938 & n13584;
  assign n15609 = n15607 & ~n15608;
  assign n15610 =  a[20]  & ~n15609;
  assign n15611 =  a[20]  & ~n15610;
  assign n15612 = ~n15609 & ~n15610;
  assign n15613 = ~n15611 & ~n15612;
  assign n15614 = n15602 & ~n15613;
  assign n15615 = ~n15600 & ~n15614;
  assign n15616 = ~n15528 & ~n15615;
  assign n15617 = ~n15525 & ~n15616;
  assign n15618 = ~n15511 & ~n15617;
  assign n15619 = n15511 & n15617;
  assign n15620 = ~n15618 & ~n15619;
  assign n15621 = n6233 & n13633;
  assign n15622 = n5663 & n13597;
  assign n15623 = n5939 & n13630;
  assign n15624 = ~n15622 & ~n15623;
  assign n15625 = ~n15621 & n15624;
  assign n15626 = n5666 & n13929;
  assign n15627 = n15625 & ~n15626;
  assign n15628 =  a[17]  & ~n15627;
  assign n15629 =  a[17]  & ~n15628;
  assign n15630 = ~n15627 & ~n15628;
  assign n15631 = ~n15629 & ~n15630;
  assign n15632 = n15620 & ~n15631;
  assign n15633 = ~n15618 & ~n15632;
  assign n15634 = ~n13438 & ~n13845;
  assign n15635 = n6402 & n13941;
  assign n15636 = ~n15634 & ~n15635;
  assign n15637 = ~n6397 & n15636;
  assign n15638 = n13951 & n15636;
  assign n15639 = ~n15637 & ~n15638;
  assign n15640 =  a[14]  & ~n15639;
  assign n15641 = ~ a[14]  & n15639;
  assign n15642 = ~n15640 & ~n15641;
  assign n15643 = ~n15633 & ~n15642;
  assign n15644 = n15472 & ~n15484;
  assign n15645 = ~n15483 & ~n15484;
  assign n15646 = ~n15644 & ~n15645;
  assign n15647 = n15633 & n15642;
  assign n15648 = ~n15643 & ~n15647;
  assign n15649 = ~n15646 & n15648;
  assign n15650 = ~n15643 & ~n15649;
  assign n15651 = ~n15499 & n15502;
  assign n15652 = ~n15503 & ~n15651;
  assign n15653 = ~n15650 & n15652;
  assign n15654 = ~n15646 & ~n15649;
  assign n15655 = n15648 & ~n15649;
  assign n15656 = ~n15654 & ~n15655;
  assign n15657 = n15620 & ~n15632;
  assign n15658 = ~n15631 & ~n15632;
  assign n15659 = ~n15657 & ~n15658;
  assign n15660 = n15528 & n15615;
  assign n15661 = ~n15616 & ~n15660;
  assign n15662 = n6233 & n13630;
  assign n15663 = n5663 & n13515;
  assign n15664 = n5939 & n13597;
  assign n15665 = ~n15663 & ~n15664;
  assign n15666 = ~n15662 & n15665;
  assign n15667 = n5666 & n13976;
  assign n15668 = n15666 & ~n15667;
  assign n15669 =  a[17]  & ~n15668;
  assign n15670 =  a[17]  & ~n15669;
  assign n15671 = ~n15668 & ~n15669;
  assign n15672 = ~n15670 & ~n15671;
  assign n15673 = n15661 & ~n15672;
  assign n15674 = n15661 & ~n15673;
  assign n15675 = ~n15672 & ~n15673;
  assign n15676 = ~n15674 & ~n15675;
  assign n15677 = n15602 & ~n15614;
  assign n15678 = ~n15613 & ~n15614;
  assign n15679 = ~n15677 & ~n15678;
  assign n15680 = n15586 & ~n15598;
  assign n15681 = ~n15597 & ~n15598;
  assign n15682 = ~n15680 & ~n15681;
  assign n15683 = n15551 & n15581;
  assign n15684 = ~n15582 & ~n15683;
  assign n15685 = n4694 & n12370;
  assign n15686 = n4533 & n12508;
  assign n15687 = n4604 & n12505;
  assign n15688 = ~n15686 & ~n15687;
  assign n15689 = ~n15685 & n15688;
  assign n15690 = n4536 & ~n13748;
  assign n15691 = n15689 & ~n15690;
  assign n15692 =  a[23]  & ~n15691;
  assign n15693 =  a[23]  & ~n15692;
  assign n15694 = ~n15691 & ~n15692;
  assign n15695 = ~n15693 & ~n15694;
  assign n15696 = n15684 & ~n15695;
  assign n15697 = n15684 & ~n15696;
  assign n15698 = ~n15695 & ~n15696;
  assign n15699 = ~n15697 & ~n15698;
  assign n15700 = ~n15568 & ~n15580;
  assign n15701 = ~n15579 & ~n15580;
  assign n15702 = ~n15700 & ~n15701;
  assign n15703 = ~n15371 & ~n15374;
  assign n15704 = ~n15372 & n15375;
  assign n15705 = ~n15703 & ~n15704;
  assign n15706 = ~n12623 & ~n12626;
  assign n15707 = ~n12624 & n12627;
  assign n15708 = ~n15706 & ~n15707;
  assign n15709 = n75 & ~n15708;
  assign n15710 = n3020 & n12540;
  assign n15711 = n3023 & n12546;
  assign n15712 = n3028 & n12543;
  assign n15713 = ~n15711 & ~n15712;
  assign n15714 = ~n15710 & n15713;
  assign n15715 = ~n15709 & n15714;
  assign n15716 = ~n15705 & ~n15715;
  assign n15717 = ~n15705 & ~n15716;
  assign n15718 = ~n15715 & ~n15716;
  assign n15719 = ~n15717 & ~n15718;
  assign n15720 = ~n15367 & ~n15370;
  assign n15721 = ~n15368 & n15371;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = n12619 & ~n12621;
  assign n15724 = ~n12622 & ~n15723;
  assign n15725 = n75 & n15724;
  assign n15726 = n3020 & n12543;
  assign n15727 = n3023 & n12549;
  assign n15728 = n3028 & n12546;
  assign n15729 = ~n15727 & ~n15728;
  assign n15730 = ~n15726 & n15729;
  assign n15731 = ~n15725 & n15730;
  assign n15732 = ~n15722 & ~n15731;
  assign n15733 = ~n15722 & ~n15732;
  assign n15734 = ~n15731 & ~n15732;
  assign n15735 = ~n15733 & ~n15734;
  assign n15736 = ~n15363 & ~n15366;
  assign n15737 = ~n15364 & n15367;
  assign n15738 = ~n15736 & ~n15737;
  assign n15739 = ~n289 & n12830;
  assign n15740 = ~n395 & n15739;
  assign n15741 = ~n173 & n15740;
  assign n15742 = ~n306 & n15741;
  assign n15743 = ~n270 & n15742;
  assign n15744 = n2784 & n3162;
  assign n15745 = n2807 & n15744;
  assign n15746 = n2262 & n15745;
  assign n15747 = n2091 & n15746;
  assign n15748 = n688 & n15747;
  assign n15749 = n4815 & n15748;
  assign n15750 = n14386 & n15749;
  assign n15751 = n15743 & n15750;
  assign n15752 = n288 & n15751;
  assign n15753 = n356 & n15752;
  assign n15754 = n116 & n15753;
  assign n15755 = ~n149 & n15754;
  assign n15756 = ~n396 & n15755;
  assign n15757 = ~n167 & n15756;
  assign n15758 = ~n99 & n15757;
  assign n15759 = ~n237 & n15758;
  assign n15760 = n3020 & n12549;
  assign n15761 = n3028 & n12552;
  assign n15762 = n3023 & n12555;
  assign n15763 = n12611 & ~n12613;
  assign n15764 = ~n12614 & ~n15763;
  assign n15765 = n75 & n15764;
  assign n15766 = ~n15762 & ~n15765;
  assign n15767 = ~n15761 & n15766;
  assign n15768 = ~n15760 & n15767;
  assign n15769 = ~n15759 & ~n15768;
  assign n15770 = n1073 & n3042;
  assign n15771 = n2704 & n15770;
  assign n15772 = n2808 & n15771;
  assign n15773 = n2422 & n15772;
  assign n15774 = n13221 & n15773;
  assign n15775 = n6026 & n15774;
  assign n15776 = n1039 & n15775;
  assign n15777 = n556 & n15776;
  assign n15778 = n230 & n15777;
  assign n15779 = n454 & n15778;
  assign n15780 = ~n301 & n15779;
  assign n15781 = ~n1101 & n15780;
  assign n15782 = ~n716 & n15781;
  assign n15783 = ~n99 & n15782;
  assign n15784 = ~n86 & n15783;
  assign n15785 = ~n429 & n15784;
  assign n15786 = n3020 & n12552;
  assign n15787 = n3028 & n12555;
  assign n15788 = n3023 & n12558;
  assign n15789 = ~n12607 & ~n12610;
  assign n15790 = ~n12608 & n12611;
  assign n15791 = ~n15789 & ~n15790;
  assign n15792 = n75 & ~n15791;
  assign n15793 = ~n15788 & ~n15792;
  assign n15794 = ~n15787 & n15793;
  assign n15795 = ~n15786 & n15794;
  assign n15796 = ~n15785 & ~n15795;
  assign n15797 = n2607 & n3987;
  assign n15798 = n1604 & n15797;
  assign n15799 = n1754 & n15798;
  assign n15800 = n2555 & n15799;
  assign n15801 = n15330 & n15800;
  assign n15802 = n874 & n15801;
  assign n15803 = n1475 & n15802;
  assign n15804 = n4295 & n15803;
  assign n15805 = n1040 & n15804;
  assign n15806 = ~n281 & n15805;
  assign n15807 = ~n641 & n15806;
  assign n15808 = ~n170 & n15807;
  assign n15809 = ~n657 & n15808;
  assign n15810 = ~n771 & n15809;
  assign n15811 = n3020 & n12555;
  assign n15812 = n3028 & n12558;
  assign n15813 = n3023 & n12561;
  assign n15814 = ~n12603 & ~n12606;
  assign n15815 = ~n12604 & n12607;
  assign n15816 = ~n15814 & ~n15815;
  assign n15817 = n75 & ~n15816;
  assign n15818 = ~n15813 & ~n15817;
  assign n15819 = ~n15812 & n15818;
  assign n15820 = ~n15811 & n15819;
  assign n15821 = ~n15810 & ~n15820;
  assign n15822 = n202 & n877;
  assign n15823 = ~n364 & n15822;
  assign n15824 = ~n339 & n15823;
  assign n15825 = ~n493 & n15824;
  assign n15826 = ~n225 & n15825;
  assign n15827 = n1272 & n1586;
  assign n15828 = n12428 & n15827;
  assign n15829 = n3219 & n15828;
  assign n15830 = n3415 & n15829;
  assign n15831 = n6769 & n15830;
  assign n15832 = n6707 & n15831;
  assign n15833 = n1916 & n15832;
  assign n15834 = n1475 & n15833;
  assign n15835 = n1531 & n15834;
  assign n15836 = n15826 & n15835;
  assign n15837 = ~n509 & n15836;
  assign n15838 = ~n352 & n15837;
  assign n15839 = ~n461 & n15838;
  assign n15840 = ~n689 & n15839;
  assign n15841 = ~n99 & n15840;
  assign n15842 = ~n277 & n15841;
  assign n15843 = n3020 & n12558;
  assign n15844 = n3028 & n12561;
  assign n15845 = n3023 & n12564;
  assign n15846 = n12599 & ~n12601;
  assign n15847 = ~n12602 & ~n15846;
  assign n15848 = n75 & n15847;
  assign n15849 = ~n15845 & ~n15848;
  assign n15850 = ~n15844 & n15849;
  assign n15851 = ~n15843 & n15850;
  assign n15852 = ~n15842 & ~n15851;
  assign n15853 = ~n374 & ~n505;
  assign n15854 = ~n1203 & n15853;
  assign n15855 = n1391 & n15854;
  assign n15856 = n690 & n15855;
  assign n15857 = n4101 & n15856;
  assign n15858 = n3159 & n15857;
  assign n15859 = n6604 & n15858;
  assign n15860 = n1522 & n15859;
  assign n15861 = ~n602 & n15860;
  assign n15862 = ~n239 & n15861;
  assign n15863 = ~n715 & n15862;
  assign n15864 = ~n167 & n15863;
  assign n15865 = ~n338 & n15864;
  assign n15866 = ~n295 & n15865;
  assign n15867 = ~n249 & n15866;
  assign n15868 = n2209 & n14518;
  assign n15869 = n4011 & n15868;
  assign n15870 = n5190 & n15869;
  assign n15871 = n6707 & n15870;
  assign n15872 = n3990 & n15871;
  assign n15873 = n2573 & n15872;
  assign n15874 = n937 & n15873;
  assign n15875 = n193 & n15874;
  assign n15876 = n570 & n15875;
  assign n15877 = ~n518 & n15876;
  assign n15878 = ~n673 & n15877;
  assign n15879 = ~n127 & n15878;
  assign n15880 = ~n358 & n15879;
  assign n15881 = ~n777 & n12711;
  assign n15882 = ~n81 & n15881;
  assign n15883 = n1274 & n2742;
  assign n15884 = n15882 & n15883;
  assign n15885 = n6517 & n15884;
  assign n15886 = n14210 & n15885;
  assign n15887 = n2703 & n15886;
  assign n15888 = n15880 & n15887;
  assign n15889 = n1915 & n15888;
  assign n15890 = n1129 & n15889;
  assign n15891 = n2583 & n15890;
  assign n15892 = n202 & n15891;
  assign n15893 = n15867 & n15892;
  assign n15894 = ~n353 & n15893;
  assign n15895 = ~n151 & n15894;
  assign n15896 = ~n495 & n15895;
  assign n15897 = ~n375 & n15896;
  assign n15898 = ~n1104 & n15897;
  assign n15899 = ~n371 & n15898;
  assign n15900 = n3020 & n12561;
  assign n15901 = n3028 & n12564;
  assign n15902 = n3023 & n12567;
  assign n15903 = ~n12595 & ~n12598;
  assign n15904 = ~n12596 & n12599;
  assign n15905 = ~n15903 & ~n15904;
  assign n15906 = n75 & ~n15905;
  assign n15907 = ~n15902 & ~n15906;
  assign n15908 = ~n15901 & n15907;
  assign n15909 = ~n15900 & n15908;
  assign n15910 = ~n15899 & ~n15909;
  assign n15911 = n12812 & n13249;
  assign n15912 = n14572 & n15911;
  assign n15913 = n247 & n15912;
  assign n15914 = n622 & n15913;
  assign n15915 = n1264 & n15914;
  assign n15916 = n1183 & n15915;
  assign n15917 = n1063 & n15916;
  assign n15918 = n1781 & n15917;
  assign n15919 = n2467 & n15918;
  assign n15920 = n634 & n15919;
  assign n15921 = ~n355 & n15920;
  assign n15922 = ~n689 & n15921;
  assign n15923 = ~n791 & n15922;
  assign n15924 = ~n394 & n15923;
  assign n15925 = n1798 & n2442;
  assign n15926 = n2022 & n15925;
  assign n15927 = n12805 & n15926;
  assign n15928 = n13041 & n15927;
  assign n15929 = n15924 & n15928;
  assign n15930 = n731 & n15929;
  assign n15931 = n978 & n15930;
  assign n15932 = ~n236 & n15931;
  assign n15933 = ~n1246 & n15932;
  assign n15934 = ~n602 & n15933;
  assign n15935 = ~n400 & n15934;
  assign n15936 = ~n192 & n15935;
  assign n15937 = ~n537 & n15936;
  assign n15938 = ~n170 & n15937;
  assign n15939 = n3020 & n12564;
  assign n15940 = n3028 & n12567;
  assign n15941 = n3023 & n12571;
  assign n15942 = ~n12592 & ~n12594;
  assign n15943 = ~n12569 & n12595;
  assign n15944 = ~n15942 & ~n15943;
  assign n15945 = n75 & ~n15944;
  assign n15946 = ~n15941 & ~n15945;
  assign n15947 = ~n15940 & n15946;
  assign n15948 = ~n15939 & n15947;
  assign n15949 = ~n15938 & ~n15948;
  assign n15950 = n3160 & n3391;
  assign n15951 = ~n1011 & n15950;
  assign n15952 = ~n168 & n15951;
  assign n15953 = ~n492 & n15952;
  assign n15954 = ~n121 & n13671;
  assign n15955 = ~n825 & n15954;
  assign n15956 = ~n173 & n15955;
  assign n15957 = n14476 & n15956;
  assign n15958 = n15953 & n15957;
  assign n15959 = n471 & n15958;
  assign n15960 = n1009 & n15959;
  assign n15961 = n2443 & n15960;
  assign n15962 = n827 & n15961;
  assign n15963 = ~n746 & n15962;
  assign n15964 = ~n154 & n15963;
  assign n15965 = ~n637 & n15964;
  assign n15966 = ~n302 & n15965;
  assign n15967 = ~n274 & n15966;
  assign n15968 = ~n466 & n15967;
  assign n15969 = ~n623 & n15968;
  assign n15970 = ~n363 & n15969;
  assign n15971 = n1388 & n2192;
  assign n15972 = n1693 & n15971;
  assign n15973 = n4819 & n15972;
  assign n15974 = n459 & n15973;
  assign n15975 = n1549 & n15974;
  assign n15976 = n2360 & n15975;
  assign n15977 = n1131 & n15976;
  assign n15978 = n15970 & n15977;
  assign n15979 = n1253 & n15978;
  assign n15980 = ~n135 & n15979;
  assign n15981 = ~n641 & n15980;
  assign n15982 = ~n417 & n15981;
  assign n15983 = ~n496 & n15982;
  assign n15984 = ~n714 & n15983;
  assign n15985 = n3020 & n12567;
  assign n15986 = n3028 & n12571;
  assign n15987 = n3023 & n12574;
  assign n15988 = n12588 & ~n12590;
  assign n15989 = ~n12591 & ~n15988;
  assign n15990 = n75 & n15989;
  assign n15991 = ~n15987 & ~n15990;
  assign n15992 = ~n15986 & n15991;
  assign n15993 = ~n15985 & n15992;
  assign n15994 = ~n15984 & ~n15993;
  assign n15995 = n2625 & n3148;
  assign n15996 = n595 & n15995;
  assign n15997 = n6565 & n15996;
  assign n15998 = n5304 & n15997;
  assign n15999 = n3205 & n15998;
  assign n16000 = n13210 & n15999;
  assign n16001 = n13135 & n16000;
  assign n16002 = n3912 & n16001;
  assign n16003 = n1916 & n16002;
  assign n16004 = n2073 & n16003;
  assign n16005 = ~n150 & n16004;
  assign n16006 = ~n563 & n16005;
  assign n16007 = ~n716 & n16006;
  assign n16008 = ~n468 & n16007;
  assign n16009 = n3020 & n12571;
  assign n16010 = n3028 & n12574;
  assign n16011 = n3023 & n12577;
  assign n16012 = n12584 & ~n12586;
  assign n16013 = ~n12587 & ~n16012;
  assign n16014 = n75 & n16013;
  assign n16015 = ~n16011 & ~n16014;
  assign n16016 = ~n16010 & n16015;
  assign n16017 = ~n16009 & n16016;
  assign n16018 = ~n16008 & ~n16017;
  assign n16019 = ~n150 & ~n713;
  assign n16020 = ~n589 & n16019;
  assign n16021 = n1409 & n16020;
  assign n16022 = n1103 & n16021;
  assign n16023 = n877 & n16022;
  assign n16024 = n808 & n16023;
  assign n16025 = n1480 & n16024;
  assign n16026 = n731 & n16025;
  assign n16027 = ~n111 & n16026;
  assign n16028 = ~n327 & n16027;
  assign n16029 = ~n430 & n16028;
  assign n16030 = ~n293 & n16029;
  assign n16031 = ~n429 & n16030;
  assign n16032 = n2992 & n12785;
  assign n16033 = n658 & n16032;
  assign n16034 = n3409 & n16033;
  assign n16035 = n16031 & n16034;
  assign n16036 = n14498 & n16035;
  assign n16037 = n15337 & n16036;
  assign n16038 = n5085 & n16037;
  assign n16039 = n1247 & n16038;
  assign n16040 = n418 & n16039;
  assign n16041 = ~n328 & n16040;
  assign n16042 = ~n511 & n16041;
  assign n16043 = ~n147 & n16042;
  assign n16044 = ~n292 & n16043;
  assign n16045 = ~n513 & n16044;
  assign n16046 = ~n395 & n16045;
  assign n16047 = ~n716 & n16046;
  assign n16048 = ~n436 & n16047;
  assign n16049 = ~n222 & n16048;
  assign n16050 = n1160 & n2191;
  assign n16051 = ~n752 & n16050;
  assign n16052 = ~n239 & n16051;
  assign n16053 = ~n146 & n16052;
  assign n16054 = ~n452 & n16053;
  assign n16055 = ~n161 & n16054;
  assign n16056 = n2007 & n3128;
  assign n16057 = n13268 & n16056;
  assign n16058 = n3905 & n16057;
  assign n16059 = n790 & n16058;
  assign n16060 = n15826 & n16059;
  assign n16061 = n16055 & n16060;
  assign n16062 = n282 & n16061;
  assign n16063 = n827 & n16062;
  assign n16064 = ~n107 & n16063;
  assign n16065 = ~n326 & n16064;
  assign n16066 = ~n81 & n16065;
  assign n16067 = ~n231 & n16066;
  assign n16068 = n1409 & n1644;
  assign n16069 = n2441 & n16068;
  assign n16070 = n2172 & n16069;
  assign n16071 = n3771 & n16070;
  assign n16072 = n2072 & n16071;
  assign n16073 = n6662 & n16072;
  assign n16074 = n2112 & n16073;
  assign n16075 = n2346 & n16074;
  assign n16076 = n16067 & n16075;
  assign n16077 = ~n746 & n16076;
  assign n16078 = ~n292 & n16077;
  assign n16079 = ~n192 & n16078;
  assign n16080 = ~n173 & n16079;
  assign n16081 = ~n436 & n16080;
  assign n16082 = n3020 & n12577;
  assign n16083 = n12577 & n12581;
  assign n16084 = ~n12577 & ~n12581;
  assign n16085 = ~n16083 & ~n16084;
  assign n16086 = n75 & ~n16085;
  assign n16087 = n3028 & ~n12581;
  assign n16088 = ~n16086 & ~n16087;
  assign n16089 = ~n16082 & n16088;
  assign n16090 = ~n16081 & ~n16089;
  assign n16091 = ~n16049 & n16090;
  assign n16092 = ~n12574 & n16083;
  assign n16093 = n12574 & ~n16083;
  assign n16094 = ~n16092 & ~n16093;
  assign n16095 = n75 & ~n16094;
  assign n16096 = n3020 & n12574;
  assign n16097 = n3023 & ~n12581;
  assign n16098 = n3028 & n12577;
  assign n16099 = ~n16097 & ~n16098;
  assign n16100 = ~n16096 & n16099;
  assign n16101 = ~n16095 & n16100;
  assign n16102 = n16049 & ~n16090;
  assign n16103 = ~n16091 & ~n16102;
  assign n16104 = ~n16101 & n16103;
  assign n16105 = ~n16091 & ~n16104;
  assign n16106 = ~n16008 & ~n16018;
  assign n16107 = ~n16017 & ~n16018;
  assign n16108 = ~n16106 & ~n16107;
  assign n16109 = ~n16105 & ~n16108;
  assign n16110 = ~n16018 & ~n16109;
  assign n16111 = ~n15984 & ~n15994;
  assign n16112 = ~n15993 & ~n15994;
  assign n16113 = ~n16111 & ~n16112;
  assign n16114 = ~n16110 & ~n16113;
  assign n16115 = ~n15994 & ~n16114;
  assign n16116 = ~n15938 & ~n15949;
  assign n16117 = ~n15948 & ~n15949;
  assign n16118 = ~n16116 & ~n16117;
  assign n16119 = ~n16115 & ~n16118;
  assign n16120 = ~n15949 & ~n16119;
  assign n16121 = ~n15899 & ~n15910;
  assign n16122 = ~n15909 & ~n15910;
  assign n16123 = ~n16121 & ~n16122;
  assign n16124 = ~n16120 & ~n16123;
  assign n16125 = ~n15910 & ~n16124;
  assign n16126 = ~n15842 & ~n15852;
  assign n16127 = ~n15851 & ~n15852;
  assign n16128 = ~n16126 & ~n16127;
  assign n16129 = ~n16125 & ~n16128;
  assign n16130 = ~n15852 & ~n16129;
  assign n16131 = ~n15810 & ~n15821;
  assign n16132 = ~n15820 & ~n15821;
  assign n16133 = ~n16131 & ~n16132;
  assign n16134 = ~n16130 & ~n16133;
  assign n16135 = ~n15821 & ~n16134;
  assign n16136 = ~n15785 & ~n15796;
  assign n16137 = ~n15795 & ~n15796;
  assign n16138 = ~n16136 & ~n16137;
  assign n16139 = ~n16135 & ~n16138;
  assign n16140 = ~n15796 & ~n16139;
  assign n16141 = ~n15759 & ~n15769;
  assign n16142 = ~n15768 & ~n15769;
  assign n16143 = ~n16141 & ~n16142;
  assign n16144 = ~n16140 & ~n16143;
  assign n16145 = ~n15769 & ~n16144;
  assign n16146 = ~n15738 & ~n16145;
  assign n16147 = n15738 & n16145;
  assign n16148 = ~n16146 & ~n16147;
  assign n16149 = n3457 & n12537;
  assign n16150 = n3542 & n12543;
  assign n16151 = n3606 & n12540;
  assign n16152 = ~n16150 & ~n16151;
  assign n16153 = ~n16149 & n16152;
  assign n16154 = ~n3368 & n16153;
  assign n16155 = n15385 & n16153;
  assign n16156 = ~n16154 & ~n16155;
  assign n16157 =  a[29]  & ~n16156;
  assign n16158 = ~ a[29]  & n16156;
  assign n16159 = ~n16157 & ~n16158;
  assign n16160 = n16148 & ~n16159;
  assign n16161 = ~n16146 & ~n16160;
  assign n16162 = ~n15735 & ~n16161;
  assign n16163 = ~n15732 & ~n16162;
  assign n16164 = ~n15719 & ~n16163;
  assign n16165 = ~n15716 & ~n16164;
  assign n16166 = n15382 & n15392;
  assign n16167 = ~n15393 & ~n16166;
  assign n16168 = ~n16165 & n16167;
  assign n16169 = n16165 & ~n16167;
  assign n16170 = ~n16168 & ~n16169;
  assign n16171 = n3457 & n12528;
  assign n16172 = n3542 & n12534;
  assign n16173 = n3606 & n12531;
  assign n16174 = ~n16172 & ~n16173;
  assign n16175 = ~n16171 & n16174;
  assign n16176 = n3368 & ~n15003;
  assign n16177 = n16175 & ~n16176;
  assign n16178 =  a[29]  & ~n16177;
  assign n16179 =  a[29]  & ~n16178;
  assign n16180 = ~n16177 & ~n16178;
  assign n16181 = ~n16179 & ~n16180;
  assign n16182 = n16170 & ~n16181;
  assign n16183 = ~n16168 & ~n16182;
  assign n16184 = ~n15400 & n15411;
  assign n16185 = ~n15412 & ~n16184;
  assign n16186 = ~n16183 & n16185;
  assign n16187 = n16183 & ~n16185;
  assign n16188 = ~n16186 & ~n16187;
  assign n16189 = n3884 & n12516;
  assign n16190 = n3967 & n12522;
  assign n16191 = n4046 & n12519;
  assign n16192 = ~n16190 & ~n16191;
  assign n16193 = ~n16189 & n16192;
  assign n16194 = n4050 & ~n14443;
  assign n16195 = n16193 & ~n16194;
  assign n16196 =  a[26]  & ~n16195;
  assign n16197 =  a[26]  & ~n16196;
  assign n16198 = ~n16195 & ~n16196;
  assign n16199 = ~n16197 & ~n16198;
  assign n16200 = n16188 & ~n16199;
  assign n16201 = ~n16186 & ~n16200;
  assign n16202 = ~n15702 & ~n16201;
  assign n16203 = n15702 & n16201;
  assign n16204 = ~n16202 & ~n16203;
  assign n16205 = n4694 & n12505;
  assign n16206 = n4533 & n12513;
  assign n16207 = n4604 & n12508;
  assign n16208 = ~n16206 & ~n16207;
  assign n16209 = ~n16205 & n16208;
  assign n16210 = n4536 & ~n14051;
  assign n16211 = n16209 & ~n16210;
  assign n16212 =  a[23]  & ~n16211;
  assign n16213 =  a[23]  & ~n16212;
  assign n16214 = ~n16211 & ~n16212;
  assign n16215 = ~n16213 & ~n16214;
  assign n16216 = n16204 & ~n16215;
  assign n16217 = ~n16202 & ~n16216;
  assign n16218 = ~n15699 & ~n16217;
  assign n16219 = ~n15696 & ~n16218;
  assign n16220 = ~n15682 & ~n16219;
  assign n16221 = n15682 & n16219;
  assign n16222 = ~n16220 & ~n16221;
  assign n16223 = n5496 & n13491;
  assign n16224 = n4935 & n12769;
  assign n16225 = n5407 & n12889;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = ~n16223 & n16226;
  assign n16228 = n4938 & ~n13503;
  assign n16229 = n16227 & ~n16228;
  assign n16230 =  a[20]  & ~n16229;
  assign n16231 =  a[20]  & ~n16230;
  assign n16232 = ~n16229 & ~n16230;
  assign n16233 = ~n16231 & ~n16232;
  assign n16234 = n16222 & ~n16233;
  assign n16235 = ~n16220 & ~n16234;
  assign n16236 = ~n15679 & ~n16235;
  assign n16237 = n15679 & n16235;
  assign n16238 = ~n16236 & ~n16237;
  assign n16239 = n6233 & n13597;
  assign n16240 = n5663 & n13521;
  assign n16241 = n5939 & n13515;
  assign n16242 = ~n16240 & ~n16241;
  assign n16243 = ~n16239 & n16242;
  assign n16244 = n5666 & ~n13612;
  assign n16245 = n16243 & ~n16244;
  assign n16246 =  a[17]  & ~n16245;
  assign n16247 =  a[17]  & ~n16246;
  assign n16248 = ~n16245 & ~n16246;
  assign n16249 = ~n16247 & ~n16248;
  assign n16250 = n16238 & ~n16249;
  assign n16251 = ~n16236 & ~n16250;
  assign n16252 = ~n15676 & ~n16251;
  assign n16253 = ~n15673 & ~n16252;
  assign n16254 = ~n15659 & ~n16253;
  assign n16255 = n15659 & n16253;
  assign n16256 = ~n16254 & ~n16255;
  assign n16257 = n7101 & ~n13438;
  assign n16258 = n6402 & ~n13627;
  assign n16259 = n6951 & n13941;
  assign n16260 = ~n16258 & ~n16259;
  assign n16261 = ~n16257 & n16260;
  assign n16262 = n6397 & n14028;
  assign n16263 = n16261 & ~n16262;
  assign n16264 =  a[14]  & ~n16263;
  assign n16265 =  a[14]  & ~n16264;
  assign n16266 = ~n16263 & ~n16264;
  assign n16267 = ~n16265 & ~n16266;
  assign n16268 = n16256 & ~n16267;
  assign n16269 = ~n16254 & ~n16268;
  assign n16270 = ~n15656 & ~n16269;
  assign n16271 = n15656 & n16269;
  assign n16272 = ~n16270 & ~n16271;
  assign n16273 = n16256 & ~n16268;
  assign n16274 = ~n16267 & ~n16268;
  assign n16275 = ~n16273 & ~n16274;
  assign n16276 = n16238 & ~n16250;
  assign n16277 = ~n16249 & ~n16250;
  assign n16278 = ~n16276 & ~n16277;
  assign n16279 = n16222 & ~n16234;
  assign n16280 = ~n16233 & ~n16234;
  assign n16281 = ~n16279 & ~n16280;
  assign n16282 = n15699 & n16217;
  assign n16283 = ~n16218 & ~n16282;
  assign n16284 = n5496 & n12889;
  assign n16285 = n4935 & n12502;
  assign n16286 = n5407 & n12769;
  assign n16287 = ~n16285 & ~n16286;
  assign n16288 = ~n16284 & n16287;
  assign n16289 = n4938 & n12895;
  assign n16290 = n16288 & ~n16289;
  assign n16291 =  a[20]  & ~n16290;
  assign n16292 =  a[20]  & ~n16291;
  assign n16293 = ~n16290 & ~n16291;
  assign n16294 = ~n16292 & ~n16293;
  assign n16295 = n16283 & ~n16294;
  assign n16296 = n16283 & ~n16295;
  assign n16297 = ~n16294 & ~n16295;
  assign n16298 = ~n16296 & ~n16297;
  assign n16299 = n16204 & ~n16216;
  assign n16300 = ~n16215 & ~n16216;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = n16188 & ~n16200;
  assign n16303 = ~n16199 & ~n16200;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = n16170 & ~n16182;
  assign n16306 = ~n16181 & ~n16182;
  assign n16307 = ~n16305 & ~n16306;
  assign n16308 = n3884 & n12519;
  assign n16309 = n3967 & n12525;
  assign n16310 = n4046 & n12522;
  assign n16311 = ~n16309 & ~n16310;
  assign n16312 = ~n16308 & n16311;
  assign n16313 = n4050 & n14454;
  assign n16314 = n16312 & ~n16313;
  assign n16315 =  a[26]  & ~n16314;
  assign n16316 =  a[26]  & ~n16315;
  assign n16317 = ~n16314 & ~n16315;
  assign n16318 = ~n16316 & ~n16317;
  assign n16319 = ~n16307 & ~n16318;
  assign n16320 = ~n16307 & ~n16319;
  assign n16321 = ~n16318 & ~n16319;
  assign n16322 = ~n16320 & ~n16321;
  assign n16323 = n15719 & n16163;
  assign n16324 = ~n16164 & ~n16323;
  assign n16325 = n3457 & n12531;
  assign n16326 = n3542 & n12537;
  assign n16327 = n3606 & n12534;
  assign n16328 = ~n16326 & ~n16327;
  assign n16329 = ~n16325 & n16328;
  assign n16330 = n3368 & n15255;
  assign n16331 = n16329 & ~n16330;
  assign n16332 =  a[29]  & ~n16331;
  assign n16333 =  a[29]  & ~n16332;
  assign n16334 = ~n16331 & ~n16332;
  assign n16335 = ~n16333 & ~n16334;
  assign n16336 = n16324 & ~n16335;
  assign n16337 = n16324 & ~n16336;
  assign n16338 = ~n16335 & ~n16336;
  assign n16339 = ~n16337 & ~n16338;
  assign n16340 = n3967 & n12528;
  assign n16341 = n4046 & n12525;
  assign n16342 = n3884 & n12522;
  assign n16343 = ~n16341 & ~n16342;
  assign n16344 = ~n16340 & n16343;
  assign n16345 = n4050 & n14837;
  assign n16346 = n16344 & ~n16345;
  assign n16347 =  a[26]  & ~n16346;
  assign n16348 =  a[26]  & ~n16347;
  assign n16349 = ~n16346 & ~n16347;
  assign n16350 = ~n16348 & ~n16349;
  assign n16351 = ~n16339 & ~n16350;
  assign n16352 = ~n16336 & ~n16351;
  assign n16353 = ~n16322 & ~n16352;
  assign n16354 = ~n16319 & ~n16353;
  assign n16355 = ~n16304 & ~n16354;
  assign n16356 = n16304 & n16354;
  assign n16357 = ~n16355 & ~n16356;
  assign n16358 = n4694 & n12508;
  assign n16359 = n4533 & n12511;
  assign n16360 = n4604 & n12513;
  assign n16361 = ~n16359 & ~n16360;
  assign n16362 = ~n16358 & n16361;
  assign n16363 = n4536 & n13863;
  assign n16364 = n16362 & ~n16363;
  assign n16365 =  a[23]  & ~n16364;
  assign n16366 =  a[23]  & ~n16365;
  assign n16367 = ~n16364 & ~n16365;
  assign n16368 = ~n16366 & ~n16367;
  assign n16369 = n16357 & ~n16368;
  assign n16370 = ~n16355 & ~n16369;
  assign n16371 = ~n16301 & ~n16370;
  assign n16372 = n16301 & n16370;
  assign n16373 = ~n16371 & ~n16372;
  assign n16374 = n5496 & n12769;
  assign n16375 = n4935 & n12370;
  assign n16376 = n5407 & n12502;
  assign n16377 = ~n16375 & ~n16376;
  assign n16378 = ~n16374 & n16377;
  assign n16379 = n4938 & n12999;
  assign n16380 = n16378 & ~n16379;
  assign n16381 =  a[20]  & ~n16380;
  assign n16382 =  a[20]  & ~n16381;
  assign n16383 = ~n16380 & ~n16381;
  assign n16384 = ~n16382 & ~n16383;
  assign n16385 = n16373 & ~n16384;
  assign n16386 = ~n16371 & ~n16385;
  assign n16387 = ~n16298 & ~n16386;
  assign n16388 = ~n16295 & ~n16387;
  assign n16389 = ~n16281 & ~n16388;
  assign n16390 = n16281 & n16388;
  assign n16391 = ~n16389 & ~n16390;
  assign n16392 = n6233 & n13515;
  assign n16393 = n5663 & n13518;
  assign n16394 = n5939 & n13521;
  assign n16395 = ~n16393 & ~n16394;
  assign n16396 = ~n16392 & n16395;
  assign n16397 = n5666 & n13541;
  assign n16398 = n16396 & ~n16397;
  assign n16399 =  a[17]  & ~n16398;
  assign n16400 =  a[17]  & ~n16399;
  assign n16401 = ~n16398 & ~n16399;
  assign n16402 = ~n16400 & ~n16401;
  assign n16403 = n16391 & ~n16402;
  assign n16404 = ~n16389 & ~n16403;
  assign n16405 = ~n16278 & ~n16404;
  assign n16406 = n16278 & n16404;
  assign n16407 = ~n16405 & ~n16406;
  assign n16408 = n7101 & ~n13627;
  assign n16409 = n6402 & n13630;
  assign n16410 = n6951 & n13633;
  assign n16411 = ~n16409 & ~n16410;
  assign n16412 = ~n16408 & n16411;
  assign n16413 = n6397 & ~n13654;
  assign n16414 = n16412 & ~n16413;
  assign n16415 =  a[14]  & ~n16414;
  assign n16416 =  a[14]  & ~n16415;
  assign n16417 = ~n16414 & ~n16415;
  assign n16418 = ~n16416 & ~n16417;
  assign n16419 = n16407 & ~n16418;
  assign n16420 = ~n16405 & ~n16419;
  assign n16421 = n7101 & n13941;
  assign n16422 = n6402 & n13633;
  assign n16423 = n6951 & ~n13627;
  assign n16424 = ~n16422 & ~n16423;
  assign n16425 = ~n16421 & n16424;
  assign n16426 = n6397 & n14136;
  assign n16427 = n16425 & ~n16426;
  assign n16428 =  a[14]  & ~n16427;
  assign n16429 =  a[14]  & ~n16428;
  assign n16430 = ~n16427 & ~n16428;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = ~n16420 & ~n16431;
  assign n16433 = n15676 & n16251;
  assign n16434 = ~n16252 & ~n16433;
  assign n16435 = ~n16420 & ~n16432;
  assign n16436 = ~n16431 & ~n16432;
  assign n16437 = ~n16435 & ~n16436;
  assign n16438 = n16434 & ~n16437;
  assign n16439 = ~n16432 & ~n16438;
  assign n16440 = ~n16275 & ~n16439;
  assign n16441 = ~n16275 & ~n16440;
  assign n16442 = ~n16439 & ~n16440;
  assign n16443 = ~n16441 & ~n16442;
  assign n16444 = n16391 & ~n16403;
  assign n16445 = ~n16402 & ~n16403;
  assign n16446 = ~n16444 & ~n16445;
  assign n16447 = n16298 & n16386;
  assign n16448 = ~n16387 & ~n16447;
  assign n16449 = n6233 & n13521;
  assign n16450 = n5663 & n13491;
  assign n16451 = n5939 & n13518;
  assign n16452 = ~n16450 & ~n16451;
  assign n16453 = ~n16449 & n16452;
  assign n16454 = n5666 & ~n13909;
  assign n16455 = n16453 & ~n16454;
  assign n16456 =  a[17]  & ~n16455;
  assign n16457 =  a[17]  & ~n16456;
  assign n16458 = ~n16455 & ~n16456;
  assign n16459 = ~n16457 & ~n16458;
  assign n16460 = n16448 & ~n16459;
  assign n16461 = n16448 & ~n16460;
  assign n16462 = ~n16459 & ~n16460;
  assign n16463 = ~n16461 & ~n16462;
  assign n16464 = n16373 & ~n16385;
  assign n16465 = ~n16384 & ~n16385;
  assign n16466 = ~n16464 & ~n16465;
  assign n16467 = n16357 & ~n16369;
  assign n16468 = ~n16368 & ~n16369;
  assign n16469 = ~n16467 & ~n16468;
  assign n16470 = n16322 & n16352;
  assign n16471 = ~n16353 & ~n16470;
  assign n16472 = n4694 & n12513;
  assign n16473 = n4533 & n12516;
  assign n16474 = n4604 & n12511;
  assign n16475 = ~n16473 & ~n16474;
  assign n16476 = ~n16472 & n16475;
  assign n16477 = n4536 & n14177;
  assign n16478 = n16476 & ~n16477;
  assign n16479 =  a[23]  & ~n16478;
  assign n16480 =  a[23]  & ~n16479;
  assign n16481 = ~n16478 & ~n16479;
  assign n16482 = ~n16480 & ~n16481;
  assign n16483 = n16471 & ~n16482;
  assign n16484 = n16471 & ~n16483;
  assign n16485 = ~n16482 & ~n16483;
  assign n16486 = ~n16484 & ~n16485;
  assign n16487 = ~n16339 & ~n16351;
  assign n16488 = ~n16350 & ~n16351;
  assign n16489 = ~n16487 & ~n16488;
  assign n16490 = n15735 & n16161;
  assign n16491 = ~n16162 & ~n16490;
  assign n16492 = n3457 & n12534;
  assign n16493 = n3542 & n12540;
  assign n16494 = n3606 & n12537;
  assign n16495 = ~n16493 & ~n16494;
  assign n16496 = ~n16492 & n16495;
  assign n16497 = n3368 & ~n15096;
  assign n16498 = n16496 & ~n16497;
  assign n16499 =  a[29]  & ~n16498;
  assign n16500 =  a[29]  & ~n16499;
  assign n16501 = ~n16498 & ~n16499;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = n16491 & ~n16502;
  assign n16504 = n16491 & ~n16503;
  assign n16505 = ~n16502 & ~n16503;
  assign n16506 = ~n16504 & ~n16505;
  assign n16507 = n4046 & n12528;
  assign n16508 = n3884 & n12525;
  assign n16509 = n3967 & n12531;
  assign n16510 = ~n16508 & ~n16509;
  assign n16511 = ~n16507 & n16510;
  assign n16512 = n4050 & n14608;
  assign n16513 = n16511 & ~n16512;
  assign n16514 =  a[26]  & ~n16513;
  assign n16515 =  a[26]  & ~n16514;
  assign n16516 = ~n16513 & ~n16514;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = ~n16506 & ~n16517;
  assign n16519 = ~n16503 & ~n16518;
  assign n16520 = ~n16489 & ~n16519;
  assign n16521 = n16489 & n16519;
  assign n16522 = ~n16520 & ~n16521;
  assign n16523 = n4694 & n12511;
  assign n16524 = n4533 & n12519;
  assign n16525 = n4604 & n12516;
  assign n16526 = ~n16524 & ~n16525;
  assign n16527 = ~n16523 & n16526;
  assign n16528 = n4536 & ~n14233;
  assign n16529 = n16527 & ~n16528;
  assign n16530 =  a[23]  & ~n16529;
  assign n16531 =  a[23]  & ~n16530;
  assign n16532 = ~n16529 & ~n16530;
  assign n16533 = ~n16531 & ~n16532;
  assign n16534 = n16522 & ~n16533;
  assign n16535 = ~n16520 & ~n16534;
  assign n16536 = ~n16486 & ~n16535;
  assign n16537 = ~n16483 & ~n16536;
  assign n16538 = ~n16469 & ~n16537;
  assign n16539 = n16469 & n16537;
  assign n16540 = ~n16538 & ~n16539;
  assign n16541 = n5496 & n12502;
  assign n16542 = n4935 & n12505;
  assign n16543 = n5407 & n12370;
  assign n16544 = ~n16542 & ~n16543;
  assign n16545 = ~n16541 & n16544;
  assign n16546 = n4938 & ~n13736;
  assign n16547 = n16545 & ~n16546;
  assign n16548 =  a[20]  & ~n16547;
  assign n16549 =  a[20]  & ~n16548;
  assign n16550 = ~n16547 & ~n16548;
  assign n16551 = ~n16549 & ~n16550;
  assign n16552 = n16540 & ~n16551;
  assign n16553 = ~n16538 & ~n16552;
  assign n16554 = ~n16466 & ~n16553;
  assign n16555 = n16466 & n16553;
  assign n16556 = ~n16554 & ~n16555;
  assign n16557 = n6233 & n13518;
  assign n16558 = n5663 & n12889;
  assign n16559 = n5939 & n13491;
  assign n16560 = ~n16558 & ~n16559;
  assign n16561 = ~n16557 & n16560;
  assign n16562 = n5666 & n13584;
  assign n16563 = n16561 & ~n16562;
  assign n16564 =  a[17]  & ~n16563;
  assign n16565 =  a[17]  & ~n16564;
  assign n16566 = ~n16563 & ~n16564;
  assign n16567 = ~n16565 & ~n16566;
  assign n16568 = n16556 & ~n16567;
  assign n16569 = ~n16554 & ~n16568;
  assign n16570 = ~n16463 & ~n16569;
  assign n16571 = ~n16460 & ~n16570;
  assign n16572 = ~n16446 & ~n16571;
  assign n16573 = n16446 & n16571;
  assign n16574 = ~n16572 & ~n16573;
  assign n16575 = n7101 & n13633;
  assign n16576 = n6402 & n13597;
  assign n16577 = n6951 & n13630;
  assign n16578 = ~n16576 & ~n16577;
  assign n16579 = ~n16575 & n16578;
  assign n16580 = n6397 & n13929;
  assign n16581 = n16579 & ~n16580;
  assign n16582 =  a[14]  & ~n16581;
  assign n16583 =  a[14]  & ~n16582;
  assign n16584 = ~n16581 & ~n16582;
  assign n16585 = ~n16583 & ~n16584;
  assign n16586 = n16574 & ~n16585;
  assign n16587 = ~n16572 & ~n16586;
  assign n16588 = ~n13438 & ~n14424;
  assign n16589 = n7291 & n13941;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = ~n7294 & n16590;
  assign n16592 = n13951 & n16590;
  assign n16593 = ~n16591 & ~n16592;
  assign n16594 =  a[11]  & ~n16593;
  assign n16595 = ~ a[11]  & n16593;
  assign n16596 = ~n16594 & ~n16595;
  assign n16597 = ~n16587 & ~n16596;
  assign n16598 = n16407 & ~n16419;
  assign n16599 = ~n16418 & ~n16419;
  assign n16600 = ~n16598 & ~n16599;
  assign n16601 = n16587 & n16596;
  assign n16602 = ~n16597 & ~n16601;
  assign n16603 = ~n16600 & n16602;
  assign n16604 = ~n16597 & ~n16603;
  assign n16605 = ~n16434 & n16437;
  assign n16606 = ~n16438 & ~n16605;
  assign n16607 = ~n16604 & n16606;
  assign n16608 = ~n16600 & ~n16603;
  assign n16609 = n16602 & ~n16603;
  assign n16610 = ~n16608 & ~n16609;
  assign n16611 = n16574 & ~n16586;
  assign n16612 = ~n16585 & ~n16586;
  assign n16613 = ~n16611 & ~n16612;
  assign n16614 = n16463 & n16569;
  assign n16615 = ~n16570 & ~n16614;
  assign n16616 = n7101 & n13630;
  assign n16617 = n6402 & n13515;
  assign n16618 = n6951 & n13597;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = ~n16616 & n16619;
  assign n16621 = n6397 & n13976;
  assign n16622 = n16620 & ~n16621;
  assign n16623 =  a[14]  & ~n16622;
  assign n16624 =  a[14]  & ~n16623;
  assign n16625 = ~n16622 & ~n16623;
  assign n16626 = ~n16624 & ~n16625;
  assign n16627 = n16615 & ~n16626;
  assign n16628 = n16615 & ~n16627;
  assign n16629 = ~n16626 & ~n16627;
  assign n16630 = ~n16628 & ~n16629;
  assign n16631 = n16556 & ~n16568;
  assign n16632 = ~n16567 & ~n16568;
  assign n16633 = ~n16631 & ~n16632;
  assign n16634 = n16540 & ~n16552;
  assign n16635 = ~n16551 & ~n16552;
  assign n16636 = ~n16634 & ~n16635;
  assign n16637 = n16486 & n16535;
  assign n16638 = ~n16536 & ~n16637;
  assign n16639 = n5496 & n12370;
  assign n16640 = n4935 & n12508;
  assign n16641 = n5407 & n12505;
  assign n16642 = ~n16640 & ~n16641;
  assign n16643 = ~n16639 & n16642;
  assign n16644 = n4938 & ~n13748;
  assign n16645 = n16643 & ~n16644;
  assign n16646 =  a[20]  & ~n16645;
  assign n16647 =  a[20]  & ~n16646;
  assign n16648 = ~n16645 & ~n16646;
  assign n16649 = ~n16647 & ~n16648;
  assign n16650 = n16638 & ~n16649;
  assign n16651 = n16638 & ~n16650;
  assign n16652 = ~n16649 & ~n16650;
  assign n16653 = ~n16651 & ~n16652;
  assign n16654 = n16522 & ~n16534;
  assign n16655 = ~n16533 & ~n16534;
  assign n16656 = ~n16654 & ~n16655;
  assign n16657 = ~n16506 & ~n16518;
  assign n16658 = ~n16517 & ~n16518;
  assign n16659 = ~n16657 & ~n16658;
  assign n16660 = ~n16140 & ~n16144;
  assign n16661 = ~n16143 & ~n16144;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = n3457 & n12540;
  assign n16664 = n3542 & n12546;
  assign n16665 = n3606 & n12543;
  assign n16666 = ~n16664 & ~n16665;
  assign n16667 = ~n16663 & n16666;
  assign n16668 = ~n3368 & n16667;
  assign n16669 = n15708 & n16667;
  assign n16670 = ~n16668 & ~n16669;
  assign n16671 =  a[29]  & ~n16670;
  assign n16672 = ~ a[29]  & n16670;
  assign n16673 = ~n16671 & ~n16672;
  assign n16674 = ~n16662 & ~n16673;
  assign n16675 = ~n16135 & ~n16139;
  assign n16676 = ~n16138 & ~n16139;
  assign n16677 = ~n16675 & ~n16676;
  assign n16678 = n3457 & n12543;
  assign n16679 = n3542 & n12549;
  assign n16680 = n3606 & n12546;
  assign n16681 = ~n16679 & ~n16680;
  assign n16682 = ~n16678 & n16681;
  assign n16683 = ~n3368 & n16682;
  assign n16684 = ~n15724 & n16682;
  assign n16685 = ~n16683 & ~n16684;
  assign n16686 =  a[29]  & ~n16685;
  assign n16687 = ~ a[29]  & n16685;
  assign n16688 = ~n16686 & ~n16687;
  assign n16689 = ~n16677 & ~n16688;
  assign n16690 = ~n16130 & ~n16134;
  assign n16691 = ~n16133 & ~n16134;
  assign n16692 = ~n16690 & ~n16691;
  assign n16693 = n3457 & n12546;
  assign n16694 = n3542 & n12552;
  assign n16695 = n3606 & n12549;
  assign n16696 = ~n16694 & ~n16695;
  assign n16697 = ~n16693 & n16696;
  assign n16698 = ~n3368 & n16697;
  assign n16699 = n15356 & n16697;
  assign n16700 = ~n16698 & ~n16699;
  assign n16701 =  a[29]  & ~n16700;
  assign n16702 = ~ a[29]  & n16700;
  assign n16703 = ~n16701 & ~n16702;
  assign n16704 = ~n16692 & ~n16703;
  assign n16705 = ~n16125 & ~n16129;
  assign n16706 = ~n16128 & ~n16129;
  assign n16707 = ~n16705 & ~n16706;
  assign n16708 = n3457 & n12549;
  assign n16709 = n3542 & n12555;
  assign n16710 = n3606 & n12552;
  assign n16711 = ~n16709 & ~n16710;
  assign n16712 = ~n16708 & n16711;
  assign n16713 = ~n3368 & n16712;
  assign n16714 = ~n15764 & n16712;
  assign n16715 = ~n16713 & ~n16714;
  assign n16716 =  a[29]  & ~n16715;
  assign n16717 = ~ a[29]  & n16715;
  assign n16718 = ~n16716 & ~n16717;
  assign n16719 = ~n16707 & ~n16718;
  assign n16720 = ~n16120 & ~n16124;
  assign n16721 = ~n16123 & ~n16124;
  assign n16722 = ~n16720 & ~n16721;
  assign n16723 = n3457 & n12552;
  assign n16724 = n3542 & n12558;
  assign n16725 = n3606 & n12555;
  assign n16726 = ~n16724 & ~n16725;
  assign n16727 = ~n16723 & n16726;
  assign n16728 = ~n3368 & n16727;
  assign n16729 = n15791 & n16727;
  assign n16730 = ~n16728 & ~n16729;
  assign n16731 =  a[29]  & ~n16730;
  assign n16732 = ~ a[29]  & n16730;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = ~n16722 & ~n16733;
  assign n16735 = n3457 & n12555;
  assign n16736 = n3542 & n12561;
  assign n16737 = n3606 & n12558;
  assign n16738 = ~n16736 & ~n16737;
  assign n16739 = ~n16735 & n16738;
  assign n16740 = n3368 & ~n15816;
  assign n16741 = n16739 & ~n16740;
  assign n16742 =  a[29]  & ~n16741;
  assign n16743 = ~n16741 & ~n16742;
  assign n16744 =  a[29]  & ~n16742;
  assign n16745 = ~n16743 & ~n16744;
  assign n16746 = ~n16115 & ~n16119;
  assign n16747 = ~n16118 & ~n16119;
  assign n16748 = ~n16746 & ~n16747;
  assign n16749 = ~n16745 & ~n16748;
  assign n16750 = ~n16745 & ~n16749;
  assign n16751 = ~n16748 & ~n16749;
  assign n16752 = ~n16750 & ~n16751;
  assign n16753 = n3457 & n12558;
  assign n16754 = n3542 & n12564;
  assign n16755 = n3606 & n12561;
  assign n16756 = ~n16754 & ~n16755;
  assign n16757 = ~n16753 & n16756;
  assign n16758 = n3368 & n15847;
  assign n16759 = n16757 & ~n16758;
  assign n16760 =  a[29]  & ~n16759;
  assign n16761 = ~n16759 & ~n16760;
  assign n16762 =  a[29]  & ~n16760;
  assign n16763 = ~n16761 & ~n16762;
  assign n16764 = ~n16110 & ~n16114;
  assign n16765 = ~n16113 & ~n16114;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = ~n16763 & ~n16766;
  assign n16768 = ~n16763 & ~n16767;
  assign n16769 = ~n16766 & ~n16767;
  assign n16770 = ~n16768 & ~n16769;
  assign n16771 = n3457 & n12561;
  assign n16772 = n3542 & n12567;
  assign n16773 = n3606 & n12564;
  assign n16774 = ~n16772 & ~n16773;
  assign n16775 = ~n16771 & n16774;
  assign n16776 = n3368 & ~n15905;
  assign n16777 = n16775 & ~n16776;
  assign n16778 =  a[29]  & ~n16777;
  assign n16779 = ~n16777 & ~n16778;
  assign n16780 =  a[29]  & ~n16778;
  assign n16781 = ~n16779 & ~n16780;
  assign n16782 = ~n16105 & ~n16109;
  assign n16783 = ~n16108 & ~n16109;
  assign n16784 = ~n16782 & ~n16783;
  assign n16785 = ~n16781 & ~n16784;
  assign n16786 = ~n16781 & ~n16785;
  assign n16787 = ~n16784 & ~n16785;
  assign n16788 = ~n16786 & ~n16787;
  assign n16789 = n3457 & n12564;
  assign n16790 = n3542 & n12571;
  assign n16791 = n3606 & n12567;
  assign n16792 = ~n16790 & ~n16791;
  assign n16793 = ~n16789 & n16792;
  assign n16794 = n3368 & ~n15944;
  assign n16795 = n16793 & ~n16794;
  assign n16796 =  a[29]  & ~n16795;
  assign n16797 = ~n16795 & ~n16796;
  assign n16798 =  a[29]  & ~n16796;
  assign n16799 = ~n16797 & ~n16798;
  assign n16800 = ~n16101 & ~n16104;
  assign n16801 = n16103 & ~n16104;
  assign n16802 = ~n16800 & ~n16801;
  assign n16803 = ~n16799 & ~n16802;
  assign n16804 = ~n16799 & ~n16803;
  assign n16805 = ~n16802 & ~n16803;
  assign n16806 = ~n16804 & ~n16805;
  assign n16807 = n3457 & n12567;
  assign n16808 = n3542 & n12574;
  assign n16809 = n3606 & n12571;
  assign n16810 = ~n16808 & ~n16809;
  assign n16811 = ~n16807 & n16810;
  assign n16812 = n3368 & n15989;
  assign n16813 = n16811 & ~n16812;
  assign n16814 =  a[29]  & ~n16813;
  assign n16815 = ~n16813 & ~n16814;
  assign n16816 =  a[29]  & ~n16814;
  assign n16817 = ~n16815 & ~n16816;
  assign n16818 = ~n16081 & ~n16090;
  assign n16819 = ~n16089 & ~n16090;
  assign n16820 = ~n16818 & ~n16819;
  assign n16821 = ~n16817 & ~n16820;
  assign n16822 = ~n16817 & ~n16821;
  assign n16823 = ~n16820 & ~n16821;
  assign n16824 = ~n16822 & ~n16823;
  assign n16825 = ~n7479 & ~n12581;
  assign n16826 = n3606 & ~n12581;
  assign n16827 = n3457 & n12577;
  assign n16828 = ~n16826 & ~n16827;
  assign n16829 = n3368 & ~n16085;
  assign n16830 = n16828 & ~n16829;
  assign n16831 =  a[29]  & ~n16830;
  assign n16832 =  a[29]  & ~n16831;
  assign n16833 = ~n16830 & ~n16831;
  assign n16834 = ~n16832 & ~n16833;
  assign n16835 = ~n3367 & ~n12581;
  assign n16836 =  a[29]  & ~n16835;
  assign n16837 = ~n16834 & n16836;
  assign n16838 = n3457 & n12574;
  assign n16839 = n3542 & ~n12581;
  assign n16840 = n3606 & n12577;
  assign n16841 = ~n16839 & ~n16840;
  assign n16842 = ~n16838 & n16841;
  assign n16843 = ~n3368 & n16842;
  assign n16844 = n16094 & n16842;
  assign n16845 = ~n16843 & ~n16844;
  assign n16846 =  a[29]  & ~n16845;
  assign n16847 = ~ a[29]  & n16845;
  assign n16848 = ~n16846 & ~n16847;
  assign n16849 = n16837 & ~n16848;
  assign n16850 = n16825 & n16849;
  assign n16851 = n3457 & n12571;
  assign n16852 = n3542 & n12577;
  assign n16853 = n3606 & n12574;
  assign n16854 = ~n16852 & ~n16853;
  assign n16855 = ~n16851 & n16854;
  assign n16856 = n3368 & n16013;
  assign n16857 = n16855 & ~n16856;
  assign n16858 =  a[29]  & ~n16857;
  assign n16859 = ~n16857 & ~n16858;
  assign n16860 =  a[29]  & ~n16858;
  assign n16861 = ~n16859 & ~n16860;
  assign n16862 = ~n16825 & n16849;
  assign n16863 = n16825 & ~n16849;
  assign n16864 = ~n16862 & ~n16863;
  assign n16865 = ~n16861 & ~n16864;
  assign n16866 = ~n16850 & ~n16865;
  assign n16867 = ~n16824 & ~n16866;
  assign n16868 = ~n16821 & ~n16867;
  assign n16869 = ~n16806 & ~n16868;
  assign n16870 = ~n16803 & ~n16869;
  assign n16871 = ~n16788 & ~n16870;
  assign n16872 = ~n16785 & ~n16871;
  assign n16873 = ~n16770 & ~n16872;
  assign n16874 = ~n16767 & ~n16873;
  assign n16875 = ~n16752 & ~n16874;
  assign n16876 = ~n16749 & ~n16875;
  assign n16877 = n16722 & n16733;
  assign n16878 = ~n16734 & ~n16877;
  assign n16879 = ~n16876 & n16878;
  assign n16880 = ~n16734 & ~n16879;
  assign n16881 = n16707 & n16718;
  assign n16882 = ~n16719 & ~n16881;
  assign n16883 = ~n16880 & n16882;
  assign n16884 = ~n16719 & ~n16883;
  assign n16885 = n16692 & n16703;
  assign n16886 = ~n16704 & ~n16885;
  assign n16887 = ~n16884 & n16886;
  assign n16888 = ~n16704 & ~n16887;
  assign n16889 = n16677 & n16688;
  assign n16890 = ~n16689 & ~n16889;
  assign n16891 = ~n16888 & n16890;
  assign n16892 = ~n16689 & ~n16891;
  assign n16893 = n16662 & n16673;
  assign n16894 = ~n16674 & ~n16893;
  assign n16895 = ~n16892 & n16894;
  assign n16896 = ~n16674 & ~n16895;
  assign n16897 = ~n16148 & n16159;
  assign n16898 = ~n16160 & ~n16897;
  assign n16899 = ~n16896 & n16898;
  assign n16900 = n16896 & ~n16898;
  assign n16901 = ~n16899 & ~n16900;
  assign n16902 = n3884 & n12528;
  assign n16903 = n3967 & n12534;
  assign n16904 = n4046 & n12531;
  assign n16905 = ~n16903 & ~n16904;
  assign n16906 = ~n16902 & n16905;
  assign n16907 = n4050 & ~n15003;
  assign n16908 = n16906 & ~n16907;
  assign n16909 =  a[26]  & ~n16908;
  assign n16910 =  a[26]  & ~n16909;
  assign n16911 = ~n16908 & ~n16909;
  assign n16912 = ~n16910 & ~n16911;
  assign n16913 = n16901 & ~n16912;
  assign n16914 = ~n16899 & ~n16913;
  assign n16915 = ~n16659 & ~n16914;
  assign n16916 = n16659 & n16914;
  assign n16917 = ~n16915 & ~n16916;
  assign n16918 = n4694 & n12516;
  assign n16919 = n4533 & n12522;
  assign n16920 = n4604 & n12519;
  assign n16921 = ~n16919 & ~n16920;
  assign n16922 = ~n16918 & n16921;
  assign n16923 = n4536 & ~n14443;
  assign n16924 = n16922 & ~n16923;
  assign n16925 =  a[23]  & ~n16924;
  assign n16926 =  a[23]  & ~n16925;
  assign n16927 = ~n16924 & ~n16925;
  assign n16928 = ~n16926 & ~n16927;
  assign n16929 = n16917 & ~n16928;
  assign n16930 = ~n16915 & ~n16929;
  assign n16931 = ~n16656 & ~n16930;
  assign n16932 = n16656 & n16930;
  assign n16933 = ~n16931 & ~n16932;
  assign n16934 = n5496 & n12505;
  assign n16935 = n4935 & n12513;
  assign n16936 = n5407 & n12508;
  assign n16937 = ~n16935 & ~n16936;
  assign n16938 = ~n16934 & n16937;
  assign n16939 = n4938 & ~n14051;
  assign n16940 = n16938 & ~n16939;
  assign n16941 =  a[20]  & ~n16940;
  assign n16942 =  a[20]  & ~n16941;
  assign n16943 = ~n16940 & ~n16941;
  assign n16944 = ~n16942 & ~n16943;
  assign n16945 = n16933 & ~n16944;
  assign n16946 = ~n16931 & ~n16945;
  assign n16947 = ~n16653 & ~n16946;
  assign n16948 = ~n16650 & ~n16947;
  assign n16949 = ~n16636 & ~n16948;
  assign n16950 = n16636 & n16948;
  assign n16951 = ~n16949 & ~n16950;
  assign n16952 = n6233 & n13491;
  assign n16953 = n5663 & n12769;
  assign n16954 = n5939 & n12889;
  assign n16955 = ~n16953 & ~n16954;
  assign n16956 = ~n16952 & n16955;
  assign n16957 = n5666 & ~n13503;
  assign n16958 = n16956 & ~n16957;
  assign n16959 =  a[17]  & ~n16958;
  assign n16960 =  a[17]  & ~n16959;
  assign n16961 = ~n16958 & ~n16959;
  assign n16962 = ~n16960 & ~n16961;
  assign n16963 = n16951 & ~n16962;
  assign n16964 = ~n16949 & ~n16963;
  assign n16965 = ~n16633 & ~n16964;
  assign n16966 = n16633 & n16964;
  assign n16967 = ~n16965 & ~n16966;
  assign n16968 = n7101 & n13597;
  assign n16969 = n6402 & n13521;
  assign n16970 = n6951 & n13515;
  assign n16971 = ~n16969 & ~n16970;
  assign n16972 = ~n16968 & n16971;
  assign n16973 = n6397 & ~n13612;
  assign n16974 = n16972 & ~n16973;
  assign n16975 =  a[14]  & ~n16974;
  assign n16976 =  a[14]  & ~n16975;
  assign n16977 = ~n16974 & ~n16975;
  assign n16978 = ~n16976 & ~n16977;
  assign n16979 = n16967 & ~n16978;
  assign n16980 = ~n16965 & ~n16979;
  assign n16981 = ~n16630 & ~n16980;
  assign n16982 = ~n16627 & ~n16981;
  assign n16983 = ~n16613 & ~n16982;
  assign n16984 = n16613 & n16982;
  assign n16985 = ~n16983 & ~n16984;
  assign n16986 = n7983 & ~n13438;
  assign n16987 = n7291 & ~n13627;
  assign n16988 = n7632 & n13941;
  assign n16989 = ~n16987 & ~n16988;
  assign n16990 = ~n16986 & n16989;
  assign n16991 = n7294 & n14028;
  assign n16992 = n16990 & ~n16991;
  assign n16993 =  a[11]  & ~n16992;
  assign n16994 =  a[11]  & ~n16993;
  assign n16995 = ~n16992 & ~n16993;
  assign n16996 = ~n16994 & ~n16995;
  assign n16997 = n16985 & ~n16996;
  assign n16998 = ~n16983 & ~n16997;
  assign n16999 = ~n16610 & ~n16998;
  assign n17000 = n16610 & n16998;
  assign n17001 = ~n16999 & ~n17000;
  assign n17002 = n16985 & ~n16997;
  assign n17003 = ~n16996 & ~n16997;
  assign n17004 = ~n17002 & ~n17003;
  assign n17005 = n16967 & ~n16979;
  assign n17006 = ~n16978 & ~n16979;
  assign n17007 = ~n17005 & ~n17006;
  assign n17008 = n16951 & ~n16963;
  assign n17009 = ~n16962 & ~n16963;
  assign n17010 = ~n17008 & ~n17009;
  assign n17011 = n16653 & n16946;
  assign n17012 = ~n16947 & ~n17011;
  assign n17013 = n6233 & n12889;
  assign n17014 = n5663 & n12502;
  assign n17015 = n5939 & n12769;
  assign n17016 = ~n17014 & ~n17015;
  assign n17017 = ~n17013 & n17016;
  assign n17018 = n5666 & n12895;
  assign n17019 = n17017 & ~n17018;
  assign n17020 =  a[17]  & ~n17019;
  assign n17021 =  a[17]  & ~n17020;
  assign n17022 = ~n17019 & ~n17020;
  assign n17023 = ~n17021 & ~n17022;
  assign n17024 = n17012 & ~n17023;
  assign n17025 = n17012 & ~n17024;
  assign n17026 = ~n17023 & ~n17024;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = n16933 & ~n16945;
  assign n17029 = ~n16944 & ~n16945;
  assign n17030 = ~n17028 & ~n17029;
  assign n17031 = n16917 & ~n16929;
  assign n17032 = ~n16928 & ~n16929;
  assign n17033 = ~n17031 & ~n17032;
  assign n17034 = n16901 & ~n16913;
  assign n17035 = ~n16912 & ~n16913;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = n16892 & ~n16894;
  assign n17038 = ~n16895 & ~n17037;
  assign n17039 = n3884 & n12531;
  assign n17040 = n3967 & n12537;
  assign n17041 = n4046 & n12534;
  assign n17042 = ~n17040 & ~n17041;
  assign n17043 = ~n17039 & n17042;
  assign n17044 = ~n4050 & n17043;
  assign n17045 = ~n15255 & n17043;
  assign n17046 = ~n17044 & ~n17045;
  assign n17047 =  a[26]  & ~n17046;
  assign n17048 = ~ a[26]  & n17046;
  assign n17049 = ~n17047 & ~n17048;
  assign n17050 = n17038 & ~n17049;
  assign n17051 = n16888 & ~n16890;
  assign n17052 = ~n16891 & ~n17051;
  assign n17053 = n3884 & n12534;
  assign n17054 = n3967 & n12540;
  assign n17055 = n4046 & n12537;
  assign n17056 = ~n17054 & ~n17055;
  assign n17057 = ~n17053 & n17056;
  assign n17058 = ~n4050 & n17057;
  assign n17059 = n15096 & n17057;
  assign n17060 = ~n17058 & ~n17059;
  assign n17061 =  a[26]  & ~n17060;
  assign n17062 = ~ a[26]  & n17060;
  assign n17063 = ~n17061 & ~n17062;
  assign n17064 = n17052 & ~n17063;
  assign n17065 = n16884 & ~n16886;
  assign n17066 = ~n16887 & ~n17065;
  assign n17067 = n3884 & n12537;
  assign n17068 = n3967 & n12543;
  assign n17069 = n4046 & n12540;
  assign n17070 = ~n17068 & ~n17069;
  assign n17071 = ~n17067 & n17070;
  assign n17072 = ~n4050 & n17071;
  assign n17073 = n15385 & n17071;
  assign n17074 = ~n17072 & ~n17073;
  assign n17075 =  a[26]  & ~n17074;
  assign n17076 = ~ a[26]  & n17074;
  assign n17077 = ~n17075 & ~n17076;
  assign n17078 = n17066 & ~n17077;
  assign n17079 = n16880 & ~n16882;
  assign n17080 = ~n16883 & ~n17079;
  assign n17081 = n3884 & n12540;
  assign n17082 = n3967 & n12546;
  assign n17083 = n4046 & n12543;
  assign n17084 = ~n17082 & ~n17083;
  assign n17085 = ~n17081 & n17084;
  assign n17086 = ~n4050 & n17085;
  assign n17087 = n15708 & n17085;
  assign n17088 = ~n17086 & ~n17087;
  assign n17089 =  a[26]  & ~n17088;
  assign n17090 = ~ a[26]  & n17088;
  assign n17091 = ~n17089 & ~n17090;
  assign n17092 = n17080 & ~n17091;
  assign n17093 = n16876 & ~n16878;
  assign n17094 = ~n16879 & ~n17093;
  assign n17095 = n3884 & n12543;
  assign n17096 = n3967 & n12549;
  assign n17097 = n4046 & n12546;
  assign n17098 = ~n17096 & ~n17097;
  assign n17099 = ~n17095 & n17098;
  assign n17100 = ~n4050 & n17099;
  assign n17101 = ~n15724 & n17099;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 =  a[26]  & ~n17102;
  assign n17104 = ~ a[26]  & n17102;
  assign n17105 = ~n17103 & ~n17104;
  assign n17106 = n17094 & ~n17105;
  assign n17107 = n16752 & n16874;
  assign n17108 = ~n16875 & ~n17107;
  assign n17109 = n3884 & n12546;
  assign n17110 = n3967 & n12552;
  assign n17111 = n4046 & n12549;
  assign n17112 = ~n17110 & ~n17111;
  assign n17113 = ~n17109 & n17112;
  assign n17114 = ~n4050 & n17113;
  assign n17115 = n15356 & n17113;
  assign n17116 = ~n17114 & ~n17115;
  assign n17117 =  a[26]  & ~n17116;
  assign n17118 = ~ a[26]  & n17116;
  assign n17119 = ~n17117 & ~n17118;
  assign n17120 = n17108 & ~n17119;
  assign n17121 = n16770 & n16872;
  assign n17122 = ~n16873 & ~n17121;
  assign n17123 = n3967 & n12555;
  assign n17124 = n4046 & n12552;
  assign n17125 = n3884 & n12549;
  assign n17126 = ~n17124 & ~n17125;
  assign n17127 = ~n17123 & n17126;
  assign n17128 = ~n4050 & n17127;
  assign n17129 = ~n15764 & n17127;
  assign n17130 = ~n17128 & ~n17129;
  assign n17131 =  a[26]  & ~n17130;
  assign n17132 = ~ a[26]  & n17130;
  assign n17133 = ~n17131 & ~n17132;
  assign n17134 = n17122 & ~n17133;
  assign n17135 = n16788 & n16870;
  assign n17136 = ~n16871 & ~n17135;
  assign n17137 = n3967 & n12558;
  assign n17138 = n3884 & n12552;
  assign n17139 = n4046 & n12555;
  assign n17140 = ~n17138 & ~n17139;
  assign n17141 = ~n17137 & n17140;
  assign n17142 = ~n4050 & n17141;
  assign n17143 = n15791 & n17141;
  assign n17144 = ~n17142 & ~n17143;
  assign n17145 =  a[26]  & ~n17144;
  assign n17146 = ~ a[26]  & n17144;
  assign n17147 = ~n17145 & ~n17146;
  assign n17148 = n17136 & ~n17147;
  assign n17149 = n16806 & n16868;
  assign n17150 = ~n16869 & ~n17149;
  assign n17151 = n4046 & n12558;
  assign n17152 = n3884 & n12555;
  assign n17153 = n3967 & n12561;
  assign n17154 = ~n17152 & ~n17153;
  assign n17155 = ~n17151 & n17154;
  assign n17156 = ~n4050 & n17155;
  assign n17157 = n15816 & n17155;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 =  a[26]  & ~n17158;
  assign n17160 = ~ a[26]  & n17158;
  assign n17161 = ~n17159 & ~n17160;
  assign n17162 = n17150 & ~n17161;
  assign n17163 = ~n16824 & ~n16867;
  assign n17164 = ~n16866 & ~n16867;
  assign n17165 = ~n17163 & ~n17164;
  assign n17166 = n3967 & n12564;
  assign n17167 = n4046 & n12561;
  assign n17168 = n3884 & n12558;
  assign n17169 = ~n17167 & ~n17168;
  assign n17170 = ~n17166 & n17169;
  assign n17171 = ~n4050 & n17170;
  assign n17172 = ~n15847 & n17170;
  assign n17173 = ~n17171 & ~n17172;
  assign n17174 =  a[26]  & ~n17173;
  assign n17175 = ~ a[26]  & n17173;
  assign n17176 = ~n17174 & ~n17175;
  assign n17177 = ~n17165 & ~n17176;
  assign n17178 = n4046 & n12564;
  assign n17179 = n3884 & n12561;
  assign n17180 = n3967 & n12567;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = ~n17178 & n17181;
  assign n17183 = n4050 & ~n15905;
  assign n17184 = n17182 & ~n17183;
  assign n17185 =  a[26]  & ~n17184;
  assign n17186 = ~n17184 & ~n17185;
  assign n17187 =  a[26]  & ~n17185;
  assign n17188 = ~n17186 & ~n17187;
  assign n17189 = n16861 & n16864;
  assign n17190 = ~n16865 & ~n17189;
  assign n17191 = ~n17188 & n17190;
  assign n17192 = ~n17188 & ~n17191;
  assign n17193 = n17190 & ~n17191;
  assign n17194 = ~n17192 & ~n17193;
  assign n17195 = n3967 & n12571;
  assign n17196 = n4046 & n12567;
  assign n17197 = n3884 & n12564;
  assign n17198 = ~n17196 & ~n17197;
  assign n17199 = ~n17195 & n17198;
  assign n17200 = n4050 & ~n15944;
  assign n17201 = n17199 & ~n17200;
  assign n17202 =  a[26]  & ~n17201;
  assign n17203 = ~n17201 & ~n17202;
  assign n17204 =  a[26]  & ~n17202;
  assign n17205 = ~n17203 & ~n17204;
  assign n17206 = ~n16837 & n16848;
  assign n17207 = ~n16849 & ~n17206;
  assign n17208 = ~n17205 & n17207;
  assign n17209 = ~n17205 & ~n17208;
  assign n17210 = n17207 & ~n17208;
  assign n17211 = ~n17209 & ~n17210;
  assign n17212 = n16834 & ~n16836;
  assign n17213 = ~n16837 & ~n17212;
  assign n17214 = n3967 & n12574;
  assign n17215 = n3884 & n12567;
  assign n17216 = n4046 & n12571;
  assign n17217 = ~n17215 & ~n17216;
  assign n17218 = ~n17214 & n17217;
  assign n17219 = ~n4050 & n17218;
  assign n17220 = ~n15989 & n17218;
  assign n17221 = ~n17219 & ~n17220;
  assign n17222 =  a[26]  & ~n17221;
  assign n17223 = ~ a[26]  & n17221;
  assign n17224 = ~n17222 & ~n17223;
  assign n17225 = n17213 & ~n17224;
  assign n17226 = n3884 & n12577;
  assign n17227 = n4046 & ~n12581;
  assign n17228 = ~n17226 & ~n17227;
  assign n17229 = n4050 & ~n16085;
  assign n17230 = n17228 & ~n17229;
  assign n17231 =  a[26]  & ~n17230;
  assign n17232 =  a[26]  & ~n17231;
  assign n17233 = ~n17230 & ~n17231;
  assign n17234 = ~n17232 & ~n17233;
  assign n17235 = ~n3880 & ~n12581;
  assign n17236 =  a[26]  & ~n17235;
  assign n17237 = ~n17234 & n17236;
  assign n17238 = n3967 & ~n12581;
  assign n17239 = n3884 & n12574;
  assign n17240 = n4046 & n12577;
  assign n17241 = ~n17239 & ~n17240;
  assign n17242 = ~n17238 & n17241;
  assign n17243 = ~n4050 & n17242;
  assign n17244 = n16094 & n17242;
  assign n17245 = ~n17243 & ~n17244;
  assign n17246 =  a[26]  & ~n17245;
  assign n17247 = ~ a[26]  & n17245;
  assign n17248 = ~n17246 & ~n17247;
  assign n17249 = n17237 & ~n17248;
  assign n17250 = n16835 & n17249;
  assign n17251 = n17249 & ~n17250;
  assign n17252 = n16835 & ~n17250;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = n3967 & n12577;
  assign n17255 = n3884 & n12571;
  assign n17256 = n4046 & n12574;
  assign n17257 = ~n17255 & ~n17256;
  assign n17258 = ~n17254 & n17257;
  assign n17259 = n4050 & n16013;
  assign n17260 = n17258 & ~n17259;
  assign n17261 =  a[26]  & ~n17260;
  assign n17262 =  a[26]  & ~n17261;
  assign n17263 = ~n17260 & ~n17261;
  assign n17264 = ~n17262 & ~n17263;
  assign n17265 = ~n17253 & ~n17264;
  assign n17266 = ~n17250 & ~n17265;
  assign n17267 = ~n17213 & n17224;
  assign n17268 = ~n17225 & ~n17267;
  assign n17269 = ~n17266 & n17268;
  assign n17270 = ~n17225 & ~n17269;
  assign n17271 = ~n17211 & ~n17270;
  assign n17272 = ~n17208 & ~n17271;
  assign n17273 = ~n17194 & ~n17272;
  assign n17274 = ~n17191 & ~n17273;
  assign n17275 = ~n17165 & ~n17177;
  assign n17276 = ~n17176 & ~n17177;
  assign n17277 = ~n17275 & ~n17276;
  assign n17278 = ~n17274 & ~n17277;
  assign n17279 = ~n17177 & ~n17278;
  assign n17280 = n17150 & ~n17162;
  assign n17281 = ~n17161 & ~n17162;
  assign n17282 = ~n17280 & ~n17281;
  assign n17283 = ~n17279 & ~n17282;
  assign n17284 = ~n17162 & ~n17283;
  assign n17285 = n17136 & ~n17148;
  assign n17286 = ~n17147 & ~n17148;
  assign n17287 = ~n17285 & ~n17286;
  assign n17288 = ~n17284 & ~n17287;
  assign n17289 = ~n17148 & ~n17288;
  assign n17290 = n17122 & ~n17134;
  assign n17291 = ~n17133 & ~n17134;
  assign n17292 = ~n17290 & ~n17291;
  assign n17293 = ~n17289 & ~n17292;
  assign n17294 = ~n17134 & ~n17293;
  assign n17295 = n17108 & ~n17120;
  assign n17296 = ~n17119 & ~n17120;
  assign n17297 = ~n17295 & ~n17296;
  assign n17298 = ~n17294 & ~n17297;
  assign n17299 = ~n17120 & ~n17298;
  assign n17300 = n17094 & ~n17106;
  assign n17301 = ~n17105 & ~n17106;
  assign n17302 = ~n17300 & ~n17301;
  assign n17303 = ~n17299 & ~n17302;
  assign n17304 = ~n17106 & ~n17303;
  assign n17305 = n17080 & ~n17092;
  assign n17306 = ~n17091 & ~n17092;
  assign n17307 = ~n17305 & ~n17306;
  assign n17308 = ~n17304 & ~n17307;
  assign n17309 = ~n17092 & ~n17308;
  assign n17310 = n17066 & ~n17078;
  assign n17311 = ~n17077 & ~n17078;
  assign n17312 = ~n17310 & ~n17311;
  assign n17313 = ~n17309 & ~n17312;
  assign n17314 = ~n17078 & ~n17313;
  assign n17315 = n17052 & ~n17064;
  assign n17316 = ~n17063 & ~n17064;
  assign n17317 = ~n17315 & ~n17316;
  assign n17318 = ~n17314 & ~n17317;
  assign n17319 = ~n17064 & ~n17318;
  assign n17320 = ~n17038 & n17049;
  assign n17321 = ~n17050 & ~n17320;
  assign n17322 = ~n17319 & n17321;
  assign n17323 = ~n17050 & ~n17322;
  assign n17324 = ~n17036 & ~n17323;
  assign n17325 = n17036 & n17323;
  assign n17326 = ~n17324 & ~n17325;
  assign n17327 = n4694 & n12519;
  assign n17328 = n4533 & n12525;
  assign n17329 = n4604 & n12522;
  assign n17330 = ~n17328 & ~n17329;
  assign n17331 = ~n17327 & n17330;
  assign n17332 = n4536 & n14454;
  assign n17333 = n17331 & ~n17332;
  assign n17334 =  a[23]  & ~n17333;
  assign n17335 =  a[23]  & ~n17334;
  assign n17336 = ~n17333 & ~n17334;
  assign n17337 = ~n17335 & ~n17336;
  assign n17338 = n17326 & ~n17337;
  assign n17339 = ~n17324 & ~n17338;
  assign n17340 = ~n17033 & ~n17339;
  assign n17341 = n17033 & n17339;
  assign n17342 = ~n17340 & ~n17341;
  assign n17343 = n5496 & n12508;
  assign n17344 = n4935 & n12511;
  assign n17345 = n5407 & n12513;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = ~n17343 & n17346;
  assign n17348 = n4938 & n13863;
  assign n17349 = n17347 & ~n17348;
  assign n17350 =  a[20]  & ~n17349;
  assign n17351 =  a[20]  & ~n17350;
  assign n17352 = ~n17349 & ~n17350;
  assign n17353 = ~n17351 & ~n17352;
  assign n17354 = n17342 & ~n17353;
  assign n17355 = ~n17340 & ~n17354;
  assign n17356 = ~n17030 & ~n17355;
  assign n17357 = n17030 & n17355;
  assign n17358 = ~n17356 & ~n17357;
  assign n17359 = n6233 & n12769;
  assign n17360 = n5663 & n12370;
  assign n17361 = n5939 & n12502;
  assign n17362 = ~n17360 & ~n17361;
  assign n17363 = ~n17359 & n17362;
  assign n17364 = n5666 & n12999;
  assign n17365 = n17363 & ~n17364;
  assign n17366 =  a[17]  & ~n17365;
  assign n17367 =  a[17]  & ~n17366;
  assign n17368 = ~n17365 & ~n17366;
  assign n17369 = ~n17367 & ~n17368;
  assign n17370 = n17358 & ~n17369;
  assign n17371 = ~n17356 & ~n17370;
  assign n17372 = ~n17027 & ~n17371;
  assign n17373 = ~n17024 & ~n17372;
  assign n17374 = ~n17010 & ~n17373;
  assign n17375 = n17010 & n17373;
  assign n17376 = ~n17374 & ~n17375;
  assign n17377 = n7101 & n13515;
  assign n17378 = n6402 & n13518;
  assign n17379 = n6951 & n13521;
  assign n17380 = ~n17378 & ~n17379;
  assign n17381 = ~n17377 & n17380;
  assign n17382 = n6397 & n13541;
  assign n17383 = n17381 & ~n17382;
  assign n17384 =  a[14]  & ~n17383;
  assign n17385 =  a[14]  & ~n17384;
  assign n17386 = ~n17383 & ~n17384;
  assign n17387 = ~n17385 & ~n17386;
  assign n17388 = n17376 & ~n17387;
  assign n17389 = ~n17374 & ~n17388;
  assign n17390 = ~n17007 & ~n17389;
  assign n17391 = n17007 & n17389;
  assign n17392 = ~n17390 & ~n17391;
  assign n17393 = n7983 & ~n13627;
  assign n17394 = n7291 & n13630;
  assign n17395 = n7632 & n13633;
  assign n17396 = ~n17394 & ~n17395;
  assign n17397 = ~n17393 & n17396;
  assign n17398 = n7294 & ~n13654;
  assign n17399 = n17397 & ~n17398;
  assign n17400 =  a[11]  & ~n17399;
  assign n17401 =  a[11]  & ~n17400;
  assign n17402 = ~n17399 & ~n17400;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = n17392 & ~n17403;
  assign n17405 = ~n17390 & ~n17404;
  assign n17406 = n7983 & n13941;
  assign n17407 = n7291 & n13633;
  assign n17408 = n7632 & ~n13627;
  assign n17409 = ~n17407 & ~n17408;
  assign n17410 = ~n17406 & n17409;
  assign n17411 = n7294 & n14136;
  assign n17412 = n17410 & ~n17411;
  assign n17413 =  a[11]  & ~n17412;
  assign n17414 =  a[11]  & ~n17413;
  assign n17415 = ~n17412 & ~n17413;
  assign n17416 = ~n17414 & ~n17415;
  assign n17417 = ~n17405 & ~n17416;
  assign n17418 = n16630 & n16980;
  assign n17419 = ~n16981 & ~n17418;
  assign n17420 = ~n17405 & ~n17417;
  assign n17421 = ~n17416 & ~n17417;
  assign n17422 = ~n17420 & ~n17421;
  assign n17423 = n17419 & ~n17422;
  assign n17424 = ~n17417 & ~n17423;
  assign n17425 = ~n17004 & ~n17424;
  assign n17426 = ~n17004 & ~n17425;
  assign n17427 = ~n17424 & ~n17425;
  assign n17428 = ~n17426 & ~n17427;
  assign n17429 = n17376 & ~n17388;
  assign n17430 = ~n17387 & ~n17388;
  assign n17431 = ~n17429 & ~n17430;
  assign n17432 = n17027 & n17371;
  assign n17433 = ~n17372 & ~n17432;
  assign n17434 = n7101 & n13521;
  assign n17435 = n6402 & n13491;
  assign n17436 = n6951 & n13518;
  assign n17437 = ~n17435 & ~n17436;
  assign n17438 = ~n17434 & n17437;
  assign n17439 = n6397 & ~n13909;
  assign n17440 = n17438 & ~n17439;
  assign n17441 =  a[14]  & ~n17440;
  assign n17442 =  a[14]  & ~n17441;
  assign n17443 = ~n17440 & ~n17441;
  assign n17444 = ~n17442 & ~n17443;
  assign n17445 = n17433 & ~n17444;
  assign n17446 = n17433 & ~n17445;
  assign n17447 = ~n17444 & ~n17445;
  assign n17448 = ~n17446 & ~n17447;
  assign n17449 = n17358 & ~n17370;
  assign n17450 = ~n17369 & ~n17370;
  assign n17451 = ~n17449 & ~n17450;
  assign n17452 = n17342 & ~n17354;
  assign n17453 = ~n17353 & ~n17354;
  assign n17454 = ~n17452 & ~n17453;
  assign n17455 = n17326 & ~n17338;
  assign n17456 = ~n17337 & ~n17338;
  assign n17457 = ~n17455 & ~n17456;
  assign n17458 = n4694 & n12522;
  assign n17459 = n4533 & n12528;
  assign n17460 = n4604 & n12525;
  assign n17461 = ~n17459 & ~n17460;
  assign n17462 = ~n17458 & n17461;
  assign n17463 = n4536 & n14837;
  assign n17464 = n17462 & ~n17463;
  assign n17465 =  a[23]  & ~n17464;
  assign n17466 = ~n17464 & ~n17465;
  assign n17467 =  a[23]  & ~n17465;
  assign n17468 = ~n17466 & ~n17467;
  assign n17469 = n17319 & ~n17321;
  assign n17470 = ~n17322 & ~n17469;
  assign n17471 = ~n17468 & n17470;
  assign n17472 = ~n17468 & ~n17471;
  assign n17473 = n17470 & ~n17471;
  assign n17474 = ~n17472 & ~n17473;
  assign n17475 = n4694 & n12525;
  assign n17476 = n4533 & n12531;
  assign n17477 = n4604 & n12528;
  assign n17478 = ~n17476 & ~n17477;
  assign n17479 = ~n17475 & n17478;
  assign n17480 = n4536 & n14608;
  assign n17481 = n17479 & ~n17480;
  assign n17482 =  a[23]  & ~n17481;
  assign n17483 = ~n17481 & ~n17482;
  assign n17484 =  a[23]  & ~n17482;
  assign n17485 = ~n17483 & ~n17484;
  assign n17486 = ~n17314 & ~n17318;
  assign n17487 = ~n17317 & ~n17318;
  assign n17488 = ~n17486 & ~n17487;
  assign n17489 = ~n17485 & ~n17488;
  assign n17490 = ~n17485 & ~n17489;
  assign n17491 = ~n17488 & ~n17489;
  assign n17492 = ~n17490 & ~n17491;
  assign n17493 = n4694 & n12528;
  assign n17494 = n4533 & n12534;
  assign n17495 = n4604 & n12531;
  assign n17496 = ~n17494 & ~n17495;
  assign n17497 = ~n17493 & n17496;
  assign n17498 = n4536 & ~n15003;
  assign n17499 = n17497 & ~n17498;
  assign n17500 =  a[23]  & ~n17499;
  assign n17501 = ~n17499 & ~n17500;
  assign n17502 =  a[23]  & ~n17500;
  assign n17503 = ~n17501 & ~n17502;
  assign n17504 = ~n17309 & ~n17313;
  assign n17505 = ~n17312 & ~n17313;
  assign n17506 = ~n17504 & ~n17505;
  assign n17507 = ~n17503 & ~n17506;
  assign n17508 = ~n17503 & ~n17507;
  assign n17509 = ~n17506 & ~n17507;
  assign n17510 = ~n17508 & ~n17509;
  assign n17511 = n4694 & n12531;
  assign n17512 = n4533 & n12537;
  assign n17513 = n4604 & n12534;
  assign n17514 = ~n17512 & ~n17513;
  assign n17515 = ~n17511 & n17514;
  assign n17516 = n4536 & n15255;
  assign n17517 = n17515 & ~n17516;
  assign n17518 =  a[23]  & ~n17517;
  assign n17519 = ~n17517 & ~n17518;
  assign n17520 =  a[23]  & ~n17518;
  assign n17521 = ~n17519 & ~n17520;
  assign n17522 = ~n17304 & ~n17308;
  assign n17523 = ~n17307 & ~n17308;
  assign n17524 = ~n17522 & ~n17523;
  assign n17525 = ~n17521 & ~n17524;
  assign n17526 = ~n17521 & ~n17525;
  assign n17527 = ~n17524 & ~n17525;
  assign n17528 = ~n17526 & ~n17527;
  assign n17529 = n4694 & n12534;
  assign n17530 = n4533 & n12540;
  assign n17531 = n4604 & n12537;
  assign n17532 = ~n17530 & ~n17531;
  assign n17533 = ~n17529 & n17532;
  assign n17534 = n4536 & ~n15096;
  assign n17535 = n17533 & ~n17534;
  assign n17536 =  a[23]  & ~n17535;
  assign n17537 = ~n17535 & ~n17536;
  assign n17538 =  a[23]  & ~n17536;
  assign n17539 = ~n17537 & ~n17538;
  assign n17540 = ~n17299 & ~n17303;
  assign n17541 = ~n17302 & ~n17303;
  assign n17542 = ~n17540 & ~n17541;
  assign n17543 = ~n17539 & ~n17542;
  assign n17544 = ~n17539 & ~n17543;
  assign n17545 = ~n17542 & ~n17543;
  assign n17546 = ~n17544 & ~n17545;
  assign n17547 = n4694 & n12537;
  assign n17548 = n4533 & n12543;
  assign n17549 = n4604 & n12540;
  assign n17550 = ~n17548 & ~n17549;
  assign n17551 = ~n17547 & n17550;
  assign n17552 = n4536 & ~n15385;
  assign n17553 = n17551 & ~n17552;
  assign n17554 =  a[23]  & ~n17553;
  assign n17555 = ~n17553 & ~n17554;
  assign n17556 =  a[23]  & ~n17554;
  assign n17557 = ~n17555 & ~n17556;
  assign n17558 = ~n17294 & ~n17298;
  assign n17559 = ~n17297 & ~n17298;
  assign n17560 = ~n17558 & ~n17559;
  assign n17561 = ~n17557 & ~n17560;
  assign n17562 = ~n17557 & ~n17561;
  assign n17563 = ~n17560 & ~n17561;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = n4694 & n12540;
  assign n17566 = n4533 & n12546;
  assign n17567 = n4604 & n12543;
  assign n17568 = ~n17566 & ~n17567;
  assign n17569 = ~n17565 & n17568;
  assign n17570 = n4536 & ~n15708;
  assign n17571 = n17569 & ~n17570;
  assign n17572 =  a[23]  & ~n17571;
  assign n17573 = ~n17571 & ~n17572;
  assign n17574 =  a[23]  & ~n17572;
  assign n17575 = ~n17573 & ~n17574;
  assign n17576 = ~n17289 & ~n17293;
  assign n17577 = ~n17292 & ~n17293;
  assign n17578 = ~n17576 & ~n17577;
  assign n17579 = ~n17575 & ~n17578;
  assign n17580 = ~n17575 & ~n17579;
  assign n17581 = ~n17578 & ~n17579;
  assign n17582 = ~n17580 & ~n17581;
  assign n17583 = n4694 & n12543;
  assign n17584 = n4533 & n12549;
  assign n17585 = n4604 & n12546;
  assign n17586 = ~n17584 & ~n17585;
  assign n17587 = ~n17583 & n17586;
  assign n17588 = n4536 & n15724;
  assign n17589 = n17587 & ~n17588;
  assign n17590 =  a[23]  & ~n17589;
  assign n17591 = ~n17589 & ~n17590;
  assign n17592 =  a[23]  & ~n17590;
  assign n17593 = ~n17591 & ~n17592;
  assign n17594 = ~n17284 & ~n17288;
  assign n17595 = ~n17287 & ~n17288;
  assign n17596 = ~n17594 & ~n17595;
  assign n17597 = ~n17593 & ~n17596;
  assign n17598 = ~n17593 & ~n17597;
  assign n17599 = ~n17596 & ~n17597;
  assign n17600 = ~n17598 & ~n17599;
  assign n17601 = n4694 & n12546;
  assign n17602 = n4533 & n12552;
  assign n17603 = n4604 & n12549;
  assign n17604 = ~n17602 & ~n17603;
  assign n17605 = ~n17601 & n17604;
  assign n17606 = n4536 & ~n15356;
  assign n17607 = n17605 & ~n17606;
  assign n17608 =  a[23]  & ~n17607;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 =  a[23]  & ~n17608;
  assign n17611 = ~n17609 & ~n17610;
  assign n17612 = ~n17279 & ~n17283;
  assign n17613 = ~n17282 & ~n17283;
  assign n17614 = ~n17612 & ~n17613;
  assign n17615 = ~n17611 & ~n17614;
  assign n17616 = ~n17611 & ~n17615;
  assign n17617 = ~n17614 & ~n17615;
  assign n17618 = ~n17616 & ~n17617;
  assign n17619 = n4694 & n12549;
  assign n17620 = n4533 & n12555;
  assign n17621 = n4604 & n12552;
  assign n17622 = ~n17620 & ~n17621;
  assign n17623 = ~n17619 & n17622;
  assign n17624 = n4536 & n15764;
  assign n17625 = n17623 & ~n17624;
  assign n17626 =  a[23]  & ~n17625;
  assign n17627 = ~n17625 & ~n17626;
  assign n17628 =  a[23]  & ~n17626;
  assign n17629 = ~n17627 & ~n17628;
  assign n17630 = ~n17274 & ~n17278;
  assign n17631 = ~n17277 & ~n17278;
  assign n17632 = ~n17630 & ~n17631;
  assign n17633 = ~n17629 & ~n17632;
  assign n17634 = ~n17629 & ~n17633;
  assign n17635 = ~n17632 & ~n17633;
  assign n17636 = ~n17634 & ~n17635;
  assign n17637 = n17194 & n17272;
  assign n17638 = ~n17273 & ~n17637;
  assign n17639 = n4694 & n12552;
  assign n17640 = n4533 & n12558;
  assign n17641 = n4604 & n12555;
  assign n17642 = ~n17640 & ~n17641;
  assign n17643 = ~n17639 & n17642;
  assign n17644 = ~n4536 & n17643;
  assign n17645 = n15791 & n17643;
  assign n17646 = ~n17644 & ~n17645;
  assign n17647 =  a[23]  & ~n17646;
  assign n17648 = ~ a[23]  & n17646;
  assign n17649 = ~n17647 & ~n17648;
  assign n17650 = n17638 & ~n17649;
  assign n17651 = n17211 & n17270;
  assign n17652 = ~n17271 & ~n17651;
  assign n17653 = n4694 & n12555;
  assign n17654 = n4533 & n12561;
  assign n17655 = n4604 & n12558;
  assign n17656 = ~n17654 & ~n17655;
  assign n17657 = ~n17653 & n17656;
  assign n17658 = ~n4536 & n17657;
  assign n17659 = n15816 & n17657;
  assign n17660 = ~n17658 & ~n17659;
  assign n17661 =  a[23]  & ~n17660;
  assign n17662 = ~ a[23]  & n17660;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = n17652 & ~n17663;
  assign n17665 = n4694 & n12558;
  assign n17666 = n4533 & n12564;
  assign n17667 = n4604 & n12561;
  assign n17668 = ~n17666 & ~n17667;
  assign n17669 = ~n17665 & n17668;
  assign n17670 = n4536 & n15847;
  assign n17671 = n17669 & ~n17670;
  assign n17672 =  a[23]  & ~n17671;
  assign n17673 = ~n17671 & ~n17672;
  assign n17674 =  a[23]  & ~n17672;
  assign n17675 = ~n17673 & ~n17674;
  assign n17676 = n17266 & ~n17268;
  assign n17677 = ~n17269 & ~n17676;
  assign n17678 = ~n17675 & n17677;
  assign n17679 = ~n17675 & ~n17678;
  assign n17680 = n17677 & ~n17678;
  assign n17681 = ~n17679 & ~n17680;
  assign n17682 = ~n17253 & ~n17265;
  assign n17683 = ~n17264 & ~n17265;
  assign n17684 = ~n17682 & ~n17683;
  assign n17685 = n4694 & n12561;
  assign n17686 = n4533 & n12567;
  assign n17687 = n4604 & n12564;
  assign n17688 = ~n17686 & ~n17687;
  assign n17689 = ~n17685 & n17688;
  assign n17690 = ~n4536 & n17689;
  assign n17691 = n15905 & n17689;
  assign n17692 = ~n17690 & ~n17691;
  assign n17693 =  a[23]  & ~n17692;
  assign n17694 = ~ a[23]  & n17692;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = ~n17684 & ~n17695;
  assign n17697 = n4694 & n12564;
  assign n17698 = n4533 & n12571;
  assign n17699 = n4604 & n12567;
  assign n17700 = ~n17698 & ~n17699;
  assign n17701 = ~n17697 & n17700;
  assign n17702 = n4536 & ~n15944;
  assign n17703 = n17701 & ~n17702;
  assign n17704 =  a[23]  & ~n17703;
  assign n17705 = ~n17703 & ~n17704;
  assign n17706 =  a[23]  & ~n17704;
  assign n17707 = ~n17705 & ~n17706;
  assign n17708 = ~n17237 & n17248;
  assign n17709 = ~n17249 & ~n17708;
  assign n17710 = ~n17707 & n17709;
  assign n17711 = ~n17707 & ~n17710;
  assign n17712 = n17709 & ~n17710;
  assign n17713 = ~n17711 & ~n17712;
  assign n17714 = n17234 & ~n17236;
  assign n17715 = ~n17237 & ~n17714;
  assign n17716 = n4694 & n12567;
  assign n17717 = n4533 & n12574;
  assign n17718 = n4604 & n12571;
  assign n17719 = ~n17717 & ~n17718;
  assign n17720 = ~n17716 & n17719;
  assign n17721 = ~n4536 & n17720;
  assign n17722 = ~n15989 & n17720;
  assign n17723 = ~n17721 & ~n17722;
  assign n17724 =  a[23]  & ~n17723;
  assign n17725 = ~ a[23]  & n17723;
  assign n17726 = ~n17724 & ~n17725;
  assign n17727 = n17715 & ~n17726;
  assign n17728 = n4604 & ~n12581;
  assign n17729 = n4694 & n12577;
  assign n17730 = ~n17728 & ~n17729;
  assign n17731 = n4536 & ~n16085;
  assign n17732 = n17730 & ~n17731;
  assign n17733 =  a[23]  & ~n17732;
  assign n17734 =  a[23]  & ~n17733;
  assign n17735 = ~n17732 & ~n17733;
  assign n17736 = ~n17734 & ~n17735;
  assign n17737 = ~n4528 & ~n12581;
  assign n17738 =  a[23]  & ~n17737;
  assign n17739 = ~n17736 & n17738;
  assign n17740 = n4694 & n12574;
  assign n17741 = n4533 & ~n12581;
  assign n17742 = n4604 & n12577;
  assign n17743 = ~n17741 & ~n17742;
  assign n17744 = ~n17740 & n17743;
  assign n17745 = ~n4536 & n17744;
  assign n17746 = n16094 & n17744;
  assign n17747 = ~n17745 & ~n17746;
  assign n17748 =  a[23]  & ~n17747;
  assign n17749 = ~ a[23]  & n17747;
  assign n17750 = ~n17748 & ~n17749;
  assign n17751 = n17739 & ~n17750;
  assign n17752 = n17235 & n17751;
  assign n17753 = n17751 & ~n17752;
  assign n17754 = n17235 & ~n17752;
  assign n17755 = ~n17753 & ~n17754;
  assign n17756 = n4694 & n12571;
  assign n17757 = n4533 & n12577;
  assign n17758 = n4604 & n12574;
  assign n17759 = ~n17757 & ~n17758;
  assign n17760 = ~n17756 & n17759;
  assign n17761 = n4536 & n16013;
  assign n17762 = n17760 & ~n17761;
  assign n17763 =  a[23]  & ~n17762;
  assign n17764 =  a[23]  & ~n17763;
  assign n17765 = ~n17762 & ~n17763;
  assign n17766 = ~n17764 & ~n17765;
  assign n17767 = ~n17755 & ~n17766;
  assign n17768 = ~n17752 & ~n17767;
  assign n17769 = ~n17715 & n17726;
  assign n17770 = ~n17727 & ~n17769;
  assign n17771 = ~n17768 & n17770;
  assign n17772 = ~n17727 & ~n17771;
  assign n17773 = ~n17713 & ~n17772;
  assign n17774 = ~n17710 & ~n17773;
  assign n17775 = n17684 & n17695;
  assign n17776 = ~n17696 & ~n17775;
  assign n17777 = ~n17774 & n17776;
  assign n17778 = ~n17696 & ~n17777;
  assign n17779 = ~n17681 & ~n17778;
  assign n17780 = ~n17678 & ~n17779;
  assign n17781 = n17652 & ~n17664;
  assign n17782 = ~n17663 & ~n17664;
  assign n17783 = ~n17781 & ~n17782;
  assign n17784 = ~n17780 & ~n17783;
  assign n17785 = ~n17664 & ~n17784;
  assign n17786 = ~n17638 & n17649;
  assign n17787 = ~n17650 & ~n17786;
  assign n17788 = ~n17785 & n17787;
  assign n17789 = ~n17650 & ~n17788;
  assign n17790 = ~n17636 & ~n17789;
  assign n17791 = ~n17633 & ~n17790;
  assign n17792 = ~n17618 & ~n17791;
  assign n17793 = ~n17615 & ~n17792;
  assign n17794 = ~n17600 & ~n17793;
  assign n17795 = ~n17597 & ~n17794;
  assign n17796 = ~n17582 & ~n17795;
  assign n17797 = ~n17579 & ~n17796;
  assign n17798 = ~n17564 & ~n17797;
  assign n17799 = ~n17561 & ~n17798;
  assign n17800 = ~n17546 & ~n17799;
  assign n17801 = ~n17543 & ~n17800;
  assign n17802 = ~n17528 & ~n17801;
  assign n17803 = ~n17525 & ~n17802;
  assign n17804 = ~n17510 & ~n17803;
  assign n17805 = ~n17507 & ~n17804;
  assign n17806 = ~n17492 & ~n17805;
  assign n17807 = ~n17489 & ~n17806;
  assign n17808 = ~n17474 & ~n17807;
  assign n17809 = ~n17471 & ~n17808;
  assign n17810 = ~n17457 & ~n17809;
  assign n17811 = n17457 & n17809;
  assign n17812 = ~n17810 & ~n17811;
  assign n17813 = n5496 & n12513;
  assign n17814 = n4935 & n12516;
  assign n17815 = n5407 & n12511;
  assign n17816 = ~n17814 & ~n17815;
  assign n17817 = ~n17813 & n17816;
  assign n17818 = n4938 & n14177;
  assign n17819 = n17817 & ~n17818;
  assign n17820 =  a[20]  & ~n17819;
  assign n17821 =  a[20]  & ~n17820;
  assign n17822 = ~n17819 & ~n17820;
  assign n17823 = ~n17821 & ~n17822;
  assign n17824 = n17812 & ~n17823;
  assign n17825 = ~n17810 & ~n17824;
  assign n17826 = ~n17454 & ~n17825;
  assign n17827 = n17454 & n17825;
  assign n17828 = ~n17826 & ~n17827;
  assign n17829 = n6233 & n12502;
  assign n17830 = n5663 & n12505;
  assign n17831 = n5939 & n12370;
  assign n17832 = ~n17830 & ~n17831;
  assign n17833 = ~n17829 & n17832;
  assign n17834 = n5666 & ~n13736;
  assign n17835 = n17833 & ~n17834;
  assign n17836 =  a[17]  & ~n17835;
  assign n17837 =  a[17]  & ~n17836;
  assign n17838 = ~n17835 & ~n17836;
  assign n17839 = ~n17837 & ~n17838;
  assign n17840 = n17828 & ~n17839;
  assign n17841 = ~n17826 & ~n17840;
  assign n17842 = ~n17451 & ~n17841;
  assign n17843 = n17451 & n17841;
  assign n17844 = ~n17842 & ~n17843;
  assign n17845 = n7101 & n13518;
  assign n17846 = n6402 & n12889;
  assign n17847 = n6951 & n13491;
  assign n17848 = ~n17846 & ~n17847;
  assign n17849 = ~n17845 & n17848;
  assign n17850 = n6397 & n13584;
  assign n17851 = n17849 & ~n17850;
  assign n17852 =  a[14]  & ~n17851;
  assign n17853 =  a[14]  & ~n17852;
  assign n17854 = ~n17851 & ~n17852;
  assign n17855 = ~n17853 & ~n17854;
  assign n17856 = n17844 & ~n17855;
  assign n17857 = ~n17842 & ~n17856;
  assign n17858 = ~n17448 & ~n17857;
  assign n17859 = ~n17445 & ~n17858;
  assign n17860 = ~n17431 & ~n17859;
  assign n17861 = n17431 & n17859;
  assign n17862 = ~n17860 & ~n17861;
  assign n17863 = n7983 & n13633;
  assign n17864 = n7291 & n13597;
  assign n17865 = n7632 & n13630;
  assign n17866 = ~n17864 & ~n17865;
  assign n17867 = ~n17863 & n17866;
  assign n17868 = n7294 & n13929;
  assign n17869 = n17867 & ~n17868;
  assign n17870 =  a[11]  & ~n17869;
  assign n17871 =  a[11]  & ~n17870;
  assign n17872 = ~n17869 & ~n17870;
  assign n17873 = ~n17871 & ~n17872;
  assign n17874 = n17862 & ~n17873;
  assign n17875 = ~n17860 & ~n17874;
  assign n17876 = ~n13438 & ~n14590;
  assign n17877 = n8418 & n13941;
  assign n17878 = ~n17876 & ~n17877;
  assign n17879 = ~n8421 & n17878;
  assign n17880 = n13951 & n17878;
  assign n17881 = ~n17879 & ~n17880;
  assign n17882 =  a[8]  & ~n17881;
  assign n17883 = ~ a[8]  & n17881;
  assign n17884 = ~n17882 & ~n17883;
  assign n17885 = ~n17875 & ~n17884;
  assign n17886 = n17392 & ~n17404;
  assign n17887 = ~n17403 & ~n17404;
  assign n17888 = ~n17886 & ~n17887;
  assign n17889 = n17875 & n17884;
  assign n17890 = ~n17885 & ~n17889;
  assign n17891 = ~n17888 & n17890;
  assign n17892 = ~n17885 & ~n17891;
  assign n17893 = ~n17419 & n17422;
  assign n17894 = ~n17423 & ~n17893;
  assign n17895 = ~n17892 & n17894;
  assign n17896 = ~n17888 & ~n17891;
  assign n17897 = n17890 & ~n17891;
  assign n17898 = ~n17896 & ~n17897;
  assign n17899 = n17862 & ~n17874;
  assign n17900 = ~n17873 & ~n17874;
  assign n17901 = ~n17899 & ~n17900;
  assign n17902 = n17448 & n17857;
  assign n17903 = ~n17858 & ~n17902;
  assign n17904 = n7983 & n13630;
  assign n17905 = n7291 & n13515;
  assign n17906 = n7632 & n13597;
  assign n17907 = ~n17905 & ~n17906;
  assign n17908 = ~n17904 & n17907;
  assign n17909 = n7294 & n13976;
  assign n17910 = n17908 & ~n17909;
  assign n17911 =  a[11]  & ~n17910;
  assign n17912 =  a[11]  & ~n17911;
  assign n17913 = ~n17910 & ~n17911;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = n17903 & ~n17914;
  assign n17916 = n17903 & ~n17915;
  assign n17917 = ~n17914 & ~n17915;
  assign n17918 = ~n17916 & ~n17917;
  assign n17919 = n17844 & ~n17856;
  assign n17920 = ~n17855 & ~n17856;
  assign n17921 = ~n17919 & ~n17920;
  assign n17922 = n17828 & ~n17840;
  assign n17923 = ~n17839 & ~n17840;
  assign n17924 = ~n17922 & ~n17923;
  assign n17925 = n17812 & ~n17824;
  assign n17926 = ~n17823 & ~n17824;
  assign n17927 = ~n17925 & ~n17926;
  assign n17928 = n17474 & n17807;
  assign n17929 = ~n17808 & ~n17928;
  assign n17930 = n5496 & n12511;
  assign n17931 = n4935 & n12519;
  assign n17932 = n5407 & n12516;
  assign n17933 = ~n17931 & ~n17932;
  assign n17934 = ~n17930 & n17933;
  assign n17935 = ~n4938 & n17934;
  assign n17936 = n14233 & n17934;
  assign n17937 = ~n17935 & ~n17936;
  assign n17938 =  a[20]  & ~n17937;
  assign n17939 = ~ a[20]  & n17937;
  assign n17940 = ~n17938 & ~n17939;
  assign n17941 = n17929 & ~n17940;
  assign n17942 = n17492 & n17805;
  assign n17943 = ~n17806 & ~n17942;
  assign n17944 = n5496 & n12516;
  assign n17945 = n4935 & n12522;
  assign n17946 = n5407 & n12519;
  assign n17947 = ~n17945 & ~n17946;
  assign n17948 = ~n17944 & n17947;
  assign n17949 = ~n4938 & n17948;
  assign n17950 = n14443 & n17948;
  assign n17951 = ~n17949 & ~n17950;
  assign n17952 =  a[20]  & ~n17951;
  assign n17953 = ~ a[20]  & n17951;
  assign n17954 = ~n17952 & ~n17953;
  assign n17955 = n17943 & ~n17954;
  assign n17956 = n17510 & n17803;
  assign n17957 = ~n17804 & ~n17956;
  assign n17958 = n5496 & n12519;
  assign n17959 = n4935 & n12525;
  assign n17960 = n5407 & n12522;
  assign n17961 = ~n17959 & ~n17960;
  assign n17962 = ~n17958 & n17961;
  assign n17963 = ~n4938 & n17962;
  assign n17964 = ~n14454 & n17962;
  assign n17965 = ~n17963 & ~n17964;
  assign n17966 =  a[20]  & ~n17965;
  assign n17967 = ~ a[20]  & n17965;
  assign n17968 = ~n17966 & ~n17967;
  assign n17969 = n17957 & ~n17968;
  assign n17970 = n17528 & n17801;
  assign n17971 = ~n17802 & ~n17970;
  assign n17972 = n5496 & n12522;
  assign n17973 = n4935 & n12528;
  assign n17974 = n5407 & n12525;
  assign n17975 = ~n17973 & ~n17974;
  assign n17976 = ~n17972 & n17975;
  assign n17977 = ~n4938 & n17976;
  assign n17978 = ~n14837 & n17976;
  assign n17979 = ~n17977 & ~n17978;
  assign n17980 =  a[20]  & ~n17979;
  assign n17981 = ~ a[20]  & n17979;
  assign n17982 = ~n17980 & ~n17981;
  assign n17983 = n17971 & ~n17982;
  assign n17984 = n17546 & n17799;
  assign n17985 = ~n17800 & ~n17984;
  assign n17986 = n5496 & n12525;
  assign n17987 = n4935 & n12531;
  assign n17988 = n5407 & n12528;
  assign n17989 = ~n17987 & ~n17988;
  assign n17990 = ~n17986 & n17989;
  assign n17991 = ~n4938 & n17990;
  assign n17992 = ~n14608 & n17990;
  assign n17993 = ~n17991 & ~n17992;
  assign n17994 =  a[20]  & ~n17993;
  assign n17995 = ~ a[20]  & n17993;
  assign n17996 = ~n17994 & ~n17995;
  assign n17997 = n17985 & ~n17996;
  assign n17998 = n17564 & n17797;
  assign n17999 = ~n17798 & ~n17998;
  assign n18000 = n5496 & n12528;
  assign n18001 = n4935 & n12534;
  assign n18002 = n5407 & n12531;
  assign n18003 = ~n18001 & ~n18002;
  assign n18004 = ~n18000 & n18003;
  assign n18005 = ~n4938 & n18004;
  assign n18006 = n15003 & n18004;
  assign n18007 = ~n18005 & ~n18006;
  assign n18008 =  a[20]  & ~n18007;
  assign n18009 = ~ a[20]  & n18007;
  assign n18010 = ~n18008 & ~n18009;
  assign n18011 = n17999 & ~n18010;
  assign n18012 = n17582 & n17795;
  assign n18013 = ~n17796 & ~n18012;
  assign n18014 = n5496 & n12531;
  assign n18015 = n4935 & n12537;
  assign n18016 = n5407 & n12534;
  assign n18017 = ~n18015 & ~n18016;
  assign n18018 = ~n18014 & n18017;
  assign n18019 = ~n4938 & n18018;
  assign n18020 = ~n15255 & n18018;
  assign n18021 = ~n18019 & ~n18020;
  assign n18022 =  a[20]  & ~n18021;
  assign n18023 = ~ a[20]  & n18021;
  assign n18024 = ~n18022 & ~n18023;
  assign n18025 = n18013 & ~n18024;
  assign n18026 = n17600 & n17793;
  assign n18027 = ~n17794 & ~n18026;
  assign n18028 = n5496 & n12534;
  assign n18029 = n4935 & n12540;
  assign n18030 = n5407 & n12537;
  assign n18031 = ~n18029 & ~n18030;
  assign n18032 = ~n18028 & n18031;
  assign n18033 = ~n4938 & n18032;
  assign n18034 = n15096 & n18032;
  assign n18035 = ~n18033 & ~n18034;
  assign n18036 =  a[20]  & ~n18035;
  assign n18037 = ~ a[20]  & n18035;
  assign n18038 = ~n18036 & ~n18037;
  assign n18039 = n18027 & ~n18038;
  assign n18040 = n17618 & n17791;
  assign n18041 = ~n17792 & ~n18040;
  assign n18042 = n5496 & n12537;
  assign n18043 = n4935 & n12543;
  assign n18044 = n5407 & n12540;
  assign n18045 = ~n18043 & ~n18044;
  assign n18046 = ~n18042 & n18045;
  assign n18047 = ~n4938 & n18046;
  assign n18048 = n15385 & n18046;
  assign n18049 = ~n18047 & ~n18048;
  assign n18050 =  a[20]  & ~n18049;
  assign n18051 = ~ a[20]  & n18049;
  assign n18052 = ~n18050 & ~n18051;
  assign n18053 = n18041 & ~n18052;
  assign n18054 = n17636 & n17789;
  assign n18055 = ~n17790 & ~n18054;
  assign n18056 = n5496 & n12540;
  assign n18057 = n4935 & n12546;
  assign n18058 = n5407 & n12543;
  assign n18059 = ~n18057 & ~n18058;
  assign n18060 = ~n18056 & n18059;
  assign n18061 = ~n4938 & n18060;
  assign n18062 = n15708 & n18060;
  assign n18063 = ~n18061 & ~n18062;
  assign n18064 =  a[20]  & ~n18063;
  assign n18065 = ~ a[20]  & n18063;
  assign n18066 = ~n18064 & ~n18065;
  assign n18067 = n18055 & ~n18066;
  assign n18068 = n5496 & n12543;
  assign n18069 = n4935 & n12549;
  assign n18070 = n5407 & n12546;
  assign n18071 = ~n18069 & ~n18070;
  assign n18072 = ~n18068 & n18071;
  assign n18073 = n4938 & n15724;
  assign n18074 = n18072 & ~n18073;
  assign n18075 =  a[20]  & ~n18074;
  assign n18076 = ~n18074 & ~n18075;
  assign n18077 =  a[20]  & ~n18075;
  assign n18078 = ~n18076 & ~n18077;
  assign n18079 = n17785 & ~n17787;
  assign n18080 = ~n17788 & ~n18079;
  assign n18081 = ~n18078 & n18080;
  assign n18082 = ~n18078 & ~n18081;
  assign n18083 = n18080 & ~n18081;
  assign n18084 = ~n18082 & ~n18083;
  assign n18085 = n5496 & n12546;
  assign n18086 = n4935 & n12552;
  assign n18087 = n5407 & n12549;
  assign n18088 = ~n18086 & ~n18087;
  assign n18089 = ~n18085 & n18088;
  assign n18090 = n4938 & ~n15356;
  assign n18091 = n18089 & ~n18090;
  assign n18092 =  a[20]  & ~n18091;
  assign n18093 = ~n18091 & ~n18092;
  assign n18094 =  a[20]  & ~n18092;
  assign n18095 = ~n18093 & ~n18094;
  assign n18096 = ~n17780 & ~n17784;
  assign n18097 = ~n17783 & ~n17784;
  assign n18098 = ~n18096 & ~n18097;
  assign n18099 = ~n18095 & ~n18098;
  assign n18100 = ~n18095 & ~n18099;
  assign n18101 = ~n18098 & ~n18099;
  assign n18102 = ~n18100 & ~n18101;
  assign n18103 = n17681 & n17778;
  assign n18104 = ~n17779 & ~n18103;
  assign n18105 = n5496 & n12549;
  assign n18106 = n4935 & n12555;
  assign n18107 = n5407 & n12552;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = ~n18105 & n18108;
  assign n18110 = ~n4938 & n18109;
  assign n18111 = ~n15764 & n18109;
  assign n18112 = ~n18110 & ~n18111;
  assign n18113 =  a[20]  & ~n18112;
  assign n18114 = ~ a[20]  & n18112;
  assign n18115 = ~n18113 & ~n18114;
  assign n18116 = n18104 & ~n18115;
  assign n18117 = n17774 & ~n17776;
  assign n18118 = ~n17777 & ~n18117;
  assign n18119 = n5496 & n12552;
  assign n18120 = n4935 & n12558;
  assign n18121 = n5407 & n12555;
  assign n18122 = ~n18120 & ~n18121;
  assign n18123 = ~n18119 & n18122;
  assign n18124 = ~n4938 & n18123;
  assign n18125 = n15791 & n18123;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 =  a[20]  & ~n18126;
  assign n18128 = ~ a[20]  & n18126;
  assign n18129 = ~n18127 & ~n18128;
  assign n18130 = n18118 & ~n18129;
  assign n18131 = n17713 & n17772;
  assign n18132 = ~n17773 & ~n18131;
  assign n18133 = n5496 & n12555;
  assign n18134 = n4935 & n12561;
  assign n18135 = n5407 & n12558;
  assign n18136 = ~n18134 & ~n18135;
  assign n18137 = ~n18133 & n18136;
  assign n18138 = ~n4938 & n18137;
  assign n18139 = n15816 & n18137;
  assign n18140 = ~n18138 & ~n18139;
  assign n18141 =  a[20]  & ~n18140;
  assign n18142 = ~ a[20]  & n18140;
  assign n18143 = ~n18141 & ~n18142;
  assign n18144 = n18132 & ~n18143;
  assign n18145 = n5496 & n12558;
  assign n18146 = n4935 & n12564;
  assign n18147 = n5407 & n12561;
  assign n18148 = ~n18146 & ~n18147;
  assign n18149 = ~n18145 & n18148;
  assign n18150 = n4938 & n15847;
  assign n18151 = n18149 & ~n18150;
  assign n18152 =  a[20]  & ~n18151;
  assign n18153 = ~n18151 & ~n18152;
  assign n18154 =  a[20]  & ~n18152;
  assign n18155 = ~n18153 & ~n18154;
  assign n18156 = n17768 & ~n17770;
  assign n18157 = ~n17771 & ~n18156;
  assign n18158 = ~n18155 & n18157;
  assign n18159 = ~n18155 & ~n18158;
  assign n18160 = n18157 & ~n18158;
  assign n18161 = ~n18159 & ~n18160;
  assign n18162 = ~n17755 & ~n17767;
  assign n18163 = ~n17766 & ~n17767;
  assign n18164 = ~n18162 & ~n18163;
  assign n18165 = n5496 & n12561;
  assign n18166 = n4935 & n12567;
  assign n18167 = n5407 & n12564;
  assign n18168 = ~n18166 & ~n18167;
  assign n18169 = ~n18165 & n18168;
  assign n18170 = ~n4938 & n18169;
  assign n18171 = n15905 & n18169;
  assign n18172 = ~n18170 & ~n18171;
  assign n18173 =  a[20]  & ~n18172;
  assign n18174 = ~ a[20]  & n18172;
  assign n18175 = ~n18173 & ~n18174;
  assign n18176 = ~n18164 & ~n18175;
  assign n18177 = n5496 & n12564;
  assign n18178 = n4935 & n12571;
  assign n18179 = n5407 & n12567;
  assign n18180 = ~n18178 & ~n18179;
  assign n18181 = ~n18177 & n18180;
  assign n18182 = n4938 & ~n15944;
  assign n18183 = n18181 & ~n18182;
  assign n18184 =  a[20]  & ~n18183;
  assign n18185 = ~n18183 & ~n18184;
  assign n18186 =  a[20]  & ~n18184;
  assign n18187 = ~n18185 & ~n18186;
  assign n18188 = ~n17739 & n17750;
  assign n18189 = ~n17751 & ~n18188;
  assign n18190 = ~n18187 & n18189;
  assign n18191 = ~n18187 & ~n18190;
  assign n18192 = n18189 & ~n18190;
  assign n18193 = ~n18191 & ~n18192;
  assign n18194 = n17736 & ~n17738;
  assign n18195 = ~n17739 & ~n18194;
  assign n18196 = n5496 & n12567;
  assign n18197 = n4935 & n12574;
  assign n18198 = n5407 & n12571;
  assign n18199 = ~n18197 & ~n18198;
  assign n18200 = ~n18196 & n18199;
  assign n18201 = ~n4938 & n18200;
  assign n18202 = ~n15989 & n18200;
  assign n18203 = ~n18201 & ~n18202;
  assign n18204 =  a[20]  & ~n18203;
  assign n18205 = ~ a[20]  & n18203;
  assign n18206 = ~n18204 & ~n18205;
  assign n18207 = n18195 & ~n18206;
  assign n18208 = n5407 & ~n12581;
  assign n18209 = n5496 & n12577;
  assign n18210 = ~n18208 & ~n18209;
  assign n18211 = n4938 & ~n16085;
  assign n18212 = n18210 & ~n18211;
  assign n18213 =  a[20]  & ~n18212;
  assign n18214 =  a[20]  & ~n18213;
  assign n18215 = ~n18212 & ~n18213;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = ~n4933 & ~n12581;
  assign n18218 =  a[20]  & ~n18217;
  assign n18219 = ~n18216 & n18218;
  assign n18220 = n5496 & n12574;
  assign n18221 = n4935 & ~n12581;
  assign n18222 = n5407 & n12577;
  assign n18223 = ~n18221 & ~n18222;
  assign n18224 = ~n18220 & n18223;
  assign n18225 = ~n4938 & n18224;
  assign n18226 = n16094 & n18224;
  assign n18227 = ~n18225 & ~n18226;
  assign n18228 =  a[20]  & ~n18227;
  assign n18229 = ~ a[20]  & n18227;
  assign n18230 = ~n18228 & ~n18229;
  assign n18231 = n18219 & ~n18230;
  assign n18232 = n17737 & n18231;
  assign n18233 = n18231 & ~n18232;
  assign n18234 = n17737 & ~n18232;
  assign n18235 = ~n18233 & ~n18234;
  assign n18236 = n5496 & n12571;
  assign n18237 = n4935 & n12577;
  assign n18238 = n5407 & n12574;
  assign n18239 = ~n18237 & ~n18238;
  assign n18240 = ~n18236 & n18239;
  assign n18241 = n4938 & n16013;
  assign n18242 = n18240 & ~n18241;
  assign n18243 =  a[20]  & ~n18242;
  assign n18244 =  a[20]  & ~n18243;
  assign n18245 = ~n18242 & ~n18243;
  assign n18246 = ~n18244 & ~n18245;
  assign n18247 = ~n18235 & ~n18246;
  assign n18248 = ~n18232 & ~n18247;
  assign n18249 = ~n18195 & n18206;
  assign n18250 = ~n18207 & ~n18249;
  assign n18251 = ~n18248 & n18250;
  assign n18252 = ~n18207 & ~n18251;
  assign n18253 = ~n18193 & ~n18252;
  assign n18254 = ~n18190 & ~n18253;
  assign n18255 = n18164 & n18175;
  assign n18256 = ~n18176 & ~n18255;
  assign n18257 = ~n18254 & n18256;
  assign n18258 = ~n18176 & ~n18257;
  assign n18259 = ~n18161 & ~n18258;
  assign n18260 = ~n18158 & ~n18259;
  assign n18261 = n18132 & ~n18144;
  assign n18262 = ~n18143 & ~n18144;
  assign n18263 = ~n18261 & ~n18262;
  assign n18264 = ~n18260 & ~n18263;
  assign n18265 = ~n18144 & ~n18264;
  assign n18266 = n18118 & ~n18130;
  assign n18267 = ~n18129 & ~n18130;
  assign n18268 = ~n18266 & ~n18267;
  assign n18269 = ~n18265 & ~n18268;
  assign n18270 = ~n18130 & ~n18269;
  assign n18271 = ~n18104 & n18115;
  assign n18272 = ~n18116 & ~n18271;
  assign n18273 = ~n18270 & n18272;
  assign n18274 = ~n18116 & ~n18273;
  assign n18275 = ~n18102 & ~n18274;
  assign n18276 = ~n18099 & ~n18275;
  assign n18277 = ~n18084 & ~n18276;
  assign n18278 = ~n18081 & ~n18277;
  assign n18279 = n18055 & ~n18067;
  assign n18280 = ~n18066 & ~n18067;
  assign n18281 = ~n18279 & ~n18280;
  assign n18282 = ~n18278 & ~n18281;
  assign n18283 = ~n18067 & ~n18282;
  assign n18284 = n18041 & ~n18053;
  assign n18285 = ~n18052 & ~n18053;
  assign n18286 = ~n18284 & ~n18285;
  assign n18287 = ~n18283 & ~n18286;
  assign n18288 = ~n18053 & ~n18287;
  assign n18289 = n18027 & ~n18039;
  assign n18290 = ~n18038 & ~n18039;
  assign n18291 = ~n18289 & ~n18290;
  assign n18292 = ~n18288 & ~n18291;
  assign n18293 = ~n18039 & ~n18292;
  assign n18294 = n18013 & ~n18025;
  assign n18295 = ~n18024 & ~n18025;
  assign n18296 = ~n18294 & ~n18295;
  assign n18297 = ~n18293 & ~n18296;
  assign n18298 = ~n18025 & ~n18297;
  assign n18299 = n17999 & ~n18011;
  assign n18300 = ~n18010 & ~n18011;
  assign n18301 = ~n18299 & ~n18300;
  assign n18302 = ~n18298 & ~n18301;
  assign n18303 = ~n18011 & ~n18302;
  assign n18304 = n17985 & ~n17997;
  assign n18305 = ~n17996 & ~n17997;
  assign n18306 = ~n18304 & ~n18305;
  assign n18307 = ~n18303 & ~n18306;
  assign n18308 = ~n17997 & ~n18307;
  assign n18309 = n17971 & ~n17983;
  assign n18310 = ~n17982 & ~n17983;
  assign n18311 = ~n18309 & ~n18310;
  assign n18312 = ~n18308 & ~n18311;
  assign n18313 = ~n17983 & ~n18312;
  assign n18314 = n17957 & ~n17969;
  assign n18315 = ~n17968 & ~n17969;
  assign n18316 = ~n18314 & ~n18315;
  assign n18317 = ~n18313 & ~n18316;
  assign n18318 = ~n17969 & ~n18317;
  assign n18319 = n17943 & ~n17955;
  assign n18320 = ~n17954 & ~n17955;
  assign n18321 = ~n18319 & ~n18320;
  assign n18322 = ~n18318 & ~n18321;
  assign n18323 = ~n17955 & ~n18322;
  assign n18324 = ~n17929 & n17940;
  assign n18325 = ~n17941 & ~n18324;
  assign n18326 = ~n18323 & n18325;
  assign n18327 = ~n17941 & ~n18326;
  assign n18328 = ~n17927 & ~n18327;
  assign n18329 = n17927 & n18327;
  assign n18330 = ~n18328 & ~n18329;
  assign n18331 = n6233 & n12370;
  assign n18332 = n5663 & n12508;
  assign n18333 = n5939 & n12505;
  assign n18334 = ~n18332 & ~n18333;
  assign n18335 = ~n18331 & n18334;
  assign n18336 = n5666 & ~n13748;
  assign n18337 = n18335 & ~n18336;
  assign n18338 =  a[17]  & ~n18337;
  assign n18339 =  a[17]  & ~n18338;
  assign n18340 = ~n18337 & ~n18338;
  assign n18341 = ~n18339 & ~n18340;
  assign n18342 = n18330 & ~n18341;
  assign n18343 = ~n18328 & ~n18342;
  assign n18344 = ~n17924 & ~n18343;
  assign n18345 = n17924 & n18343;
  assign n18346 = ~n18344 & ~n18345;
  assign n18347 = n7101 & n13491;
  assign n18348 = n6402 & n12769;
  assign n18349 = n6951 & n12889;
  assign n18350 = ~n18348 & ~n18349;
  assign n18351 = ~n18347 & n18350;
  assign n18352 = n6397 & ~n13503;
  assign n18353 = n18351 & ~n18352;
  assign n18354 =  a[14]  & ~n18353;
  assign n18355 =  a[14]  & ~n18354;
  assign n18356 = ~n18353 & ~n18354;
  assign n18357 = ~n18355 & ~n18356;
  assign n18358 = n18346 & ~n18357;
  assign n18359 = ~n18344 & ~n18358;
  assign n18360 = ~n17921 & ~n18359;
  assign n18361 = n17921 & n18359;
  assign n18362 = ~n18360 & ~n18361;
  assign n18363 = n7983 & n13597;
  assign n18364 = n7291 & n13521;
  assign n18365 = n7632 & n13515;
  assign n18366 = ~n18364 & ~n18365;
  assign n18367 = ~n18363 & n18366;
  assign n18368 = n7294 & ~n13612;
  assign n18369 = n18367 & ~n18368;
  assign n18370 =  a[11]  & ~n18369;
  assign n18371 =  a[11]  & ~n18370;
  assign n18372 = ~n18369 & ~n18370;
  assign n18373 = ~n18371 & ~n18372;
  assign n18374 = n18362 & ~n18373;
  assign n18375 = ~n18360 & ~n18374;
  assign n18376 = ~n17918 & ~n18375;
  assign n18377 = ~n17915 & ~n18376;
  assign n18378 = ~n17901 & ~n18377;
  assign n18379 = n17901 & n18377;
  assign n18380 = ~n18378 & ~n18379;
  assign n18381 = n9331 & ~n13438;
  assign n18382 = n8418 & ~n13627;
  assign n18383 = n8860 & n13941;
  assign n18384 = ~n18382 & ~n18383;
  assign n18385 = ~n18381 & n18384;
  assign n18386 = n8421 & n14028;
  assign n18387 = n18385 & ~n18386;
  assign n18388 =  a[8]  & ~n18387;
  assign n18389 =  a[8]  & ~n18388;
  assign n18390 = ~n18387 & ~n18388;
  assign n18391 = ~n18389 & ~n18390;
  assign n18392 = n18380 & ~n18391;
  assign n18393 = ~n18378 & ~n18392;
  assign n18394 = ~n17898 & ~n18393;
  assign n18395 = n17898 & n18393;
  assign n18396 = ~n18394 & ~n18395;
  assign n18397 = n18380 & ~n18392;
  assign n18398 = ~n18391 & ~n18392;
  assign n18399 = ~n18397 & ~n18398;
  assign n18400 = n18362 & ~n18374;
  assign n18401 = ~n18373 & ~n18374;
  assign n18402 = ~n18400 & ~n18401;
  assign n18403 = n18346 & ~n18358;
  assign n18404 = ~n18357 & ~n18358;
  assign n18405 = ~n18403 & ~n18404;
  assign n18406 = n18330 & ~n18342;
  assign n18407 = ~n18341 & ~n18342;
  assign n18408 = ~n18406 & ~n18407;
  assign n18409 = n6233 & n12505;
  assign n18410 = n5663 & n12513;
  assign n18411 = n5939 & n12508;
  assign n18412 = ~n18410 & ~n18411;
  assign n18413 = ~n18409 & n18412;
  assign n18414 = n5666 & ~n14051;
  assign n18415 = n18413 & ~n18414;
  assign n18416 =  a[17]  & ~n18415;
  assign n18417 = ~n18415 & ~n18416;
  assign n18418 =  a[17]  & ~n18416;
  assign n18419 = ~n18417 & ~n18418;
  assign n18420 = n18323 & ~n18325;
  assign n18421 = ~n18326 & ~n18420;
  assign n18422 = ~n18419 & n18421;
  assign n18423 = ~n18419 & ~n18422;
  assign n18424 = n18421 & ~n18422;
  assign n18425 = ~n18423 & ~n18424;
  assign n18426 = n6233 & n12508;
  assign n18427 = n5663 & n12511;
  assign n18428 = n5939 & n12513;
  assign n18429 = ~n18427 & ~n18428;
  assign n18430 = ~n18426 & n18429;
  assign n18431 = n5666 & n13863;
  assign n18432 = n18430 & ~n18431;
  assign n18433 =  a[17]  & ~n18432;
  assign n18434 = ~n18432 & ~n18433;
  assign n18435 =  a[17]  & ~n18433;
  assign n18436 = ~n18434 & ~n18435;
  assign n18437 = ~n18318 & ~n18322;
  assign n18438 = ~n18321 & ~n18322;
  assign n18439 = ~n18437 & ~n18438;
  assign n18440 = ~n18436 & ~n18439;
  assign n18441 = ~n18436 & ~n18440;
  assign n18442 = ~n18439 & ~n18440;
  assign n18443 = ~n18441 & ~n18442;
  assign n18444 = n6233 & n12513;
  assign n18445 = n5663 & n12516;
  assign n18446 = n5939 & n12511;
  assign n18447 = ~n18445 & ~n18446;
  assign n18448 = ~n18444 & n18447;
  assign n18449 = n5666 & n14177;
  assign n18450 = n18448 & ~n18449;
  assign n18451 =  a[17]  & ~n18450;
  assign n18452 = ~n18450 & ~n18451;
  assign n18453 =  a[17]  & ~n18451;
  assign n18454 = ~n18452 & ~n18453;
  assign n18455 = ~n18313 & ~n18317;
  assign n18456 = ~n18316 & ~n18317;
  assign n18457 = ~n18455 & ~n18456;
  assign n18458 = ~n18454 & ~n18457;
  assign n18459 = ~n18454 & ~n18458;
  assign n18460 = ~n18457 & ~n18458;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = n6233 & n12511;
  assign n18463 = n5663 & n12519;
  assign n18464 = n5939 & n12516;
  assign n18465 = ~n18463 & ~n18464;
  assign n18466 = ~n18462 & n18465;
  assign n18467 = n5666 & ~n14233;
  assign n18468 = n18466 & ~n18467;
  assign n18469 =  a[17]  & ~n18468;
  assign n18470 = ~n18468 & ~n18469;
  assign n18471 =  a[17]  & ~n18469;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = ~n18308 & ~n18312;
  assign n18474 = ~n18311 & ~n18312;
  assign n18475 = ~n18473 & ~n18474;
  assign n18476 = ~n18472 & ~n18475;
  assign n18477 = ~n18472 & ~n18476;
  assign n18478 = ~n18475 & ~n18476;
  assign n18479 = ~n18477 & ~n18478;
  assign n18480 = n6233 & n12516;
  assign n18481 = n5663 & n12522;
  assign n18482 = n5939 & n12519;
  assign n18483 = ~n18481 & ~n18482;
  assign n18484 = ~n18480 & n18483;
  assign n18485 = n5666 & ~n14443;
  assign n18486 = n18484 & ~n18485;
  assign n18487 =  a[17]  & ~n18486;
  assign n18488 = ~n18486 & ~n18487;
  assign n18489 =  a[17]  & ~n18487;
  assign n18490 = ~n18488 & ~n18489;
  assign n18491 = ~n18303 & ~n18307;
  assign n18492 = ~n18306 & ~n18307;
  assign n18493 = ~n18491 & ~n18492;
  assign n18494 = ~n18490 & ~n18493;
  assign n18495 = ~n18490 & ~n18494;
  assign n18496 = ~n18493 & ~n18494;
  assign n18497 = ~n18495 & ~n18496;
  assign n18498 = n6233 & n12519;
  assign n18499 = n5663 & n12525;
  assign n18500 = n5939 & n12522;
  assign n18501 = ~n18499 & ~n18500;
  assign n18502 = ~n18498 & n18501;
  assign n18503 = n5666 & n14454;
  assign n18504 = n18502 & ~n18503;
  assign n18505 =  a[17]  & ~n18504;
  assign n18506 = ~n18504 & ~n18505;
  assign n18507 =  a[17]  & ~n18505;
  assign n18508 = ~n18506 & ~n18507;
  assign n18509 = ~n18298 & ~n18302;
  assign n18510 = ~n18301 & ~n18302;
  assign n18511 = ~n18509 & ~n18510;
  assign n18512 = ~n18508 & ~n18511;
  assign n18513 = ~n18508 & ~n18512;
  assign n18514 = ~n18511 & ~n18512;
  assign n18515 = ~n18513 & ~n18514;
  assign n18516 = n6233 & n12522;
  assign n18517 = n5663 & n12528;
  assign n18518 = n5939 & n12525;
  assign n18519 = ~n18517 & ~n18518;
  assign n18520 = ~n18516 & n18519;
  assign n18521 = n5666 & n14837;
  assign n18522 = n18520 & ~n18521;
  assign n18523 =  a[17]  & ~n18522;
  assign n18524 = ~n18522 & ~n18523;
  assign n18525 =  a[17]  & ~n18523;
  assign n18526 = ~n18524 & ~n18525;
  assign n18527 = ~n18293 & ~n18297;
  assign n18528 = ~n18296 & ~n18297;
  assign n18529 = ~n18527 & ~n18528;
  assign n18530 = ~n18526 & ~n18529;
  assign n18531 = ~n18526 & ~n18530;
  assign n18532 = ~n18529 & ~n18530;
  assign n18533 = ~n18531 & ~n18532;
  assign n18534 = n6233 & n12525;
  assign n18535 = n5663 & n12531;
  assign n18536 = n5939 & n12528;
  assign n18537 = ~n18535 & ~n18536;
  assign n18538 = ~n18534 & n18537;
  assign n18539 = n5666 & n14608;
  assign n18540 = n18538 & ~n18539;
  assign n18541 =  a[17]  & ~n18540;
  assign n18542 = ~n18540 & ~n18541;
  assign n18543 =  a[17]  & ~n18541;
  assign n18544 = ~n18542 & ~n18543;
  assign n18545 = ~n18288 & ~n18292;
  assign n18546 = ~n18291 & ~n18292;
  assign n18547 = ~n18545 & ~n18546;
  assign n18548 = ~n18544 & ~n18547;
  assign n18549 = ~n18544 & ~n18548;
  assign n18550 = ~n18547 & ~n18548;
  assign n18551 = ~n18549 & ~n18550;
  assign n18552 = n6233 & n12528;
  assign n18553 = n5663 & n12534;
  assign n18554 = n5939 & n12531;
  assign n18555 = ~n18553 & ~n18554;
  assign n18556 = ~n18552 & n18555;
  assign n18557 = n5666 & ~n15003;
  assign n18558 = n18556 & ~n18557;
  assign n18559 =  a[17]  & ~n18558;
  assign n18560 = ~n18558 & ~n18559;
  assign n18561 =  a[17]  & ~n18559;
  assign n18562 = ~n18560 & ~n18561;
  assign n18563 = ~n18283 & ~n18287;
  assign n18564 = ~n18286 & ~n18287;
  assign n18565 = ~n18563 & ~n18564;
  assign n18566 = ~n18562 & ~n18565;
  assign n18567 = ~n18562 & ~n18566;
  assign n18568 = ~n18565 & ~n18566;
  assign n18569 = ~n18567 & ~n18568;
  assign n18570 = n6233 & n12531;
  assign n18571 = n5663 & n12537;
  assign n18572 = n5939 & n12534;
  assign n18573 = ~n18571 & ~n18572;
  assign n18574 = ~n18570 & n18573;
  assign n18575 = n5666 & n15255;
  assign n18576 = n18574 & ~n18575;
  assign n18577 =  a[17]  & ~n18576;
  assign n18578 = ~n18576 & ~n18577;
  assign n18579 =  a[17]  & ~n18577;
  assign n18580 = ~n18578 & ~n18579;
  assign n18581 = ~n18278 & ~n18282;
  assign n18582 = ~n18281 & ~n18282;
  assign n18583 = ~n18581 & ~n18582;
  assign n18584 = ~n18580 & ~n18583;
  assign n18585 = ~n18580 & ~n18584;
  assign n18586 = ~n18583 & ~n18584;
  assign n18587 = ~n18585 & ~n18586;
  assign n18588 = n18084 & n18276;
  assign n18589 = ~n18277 & ~n18588;
  assign n18590 = n6233 & n12534;
  assign n18591 = n5663 & n12540;
  assign n18592 = n5939 & n12537;
  assign n18593 = ~n18591 & ~n18592;
  assign n18594 = ~n18590 & n18593;
  assign n18595 = ~n5666 & n18594;
  assign n18596 = n15096 & n18594;
  assign n18597 = ~n18595 & ~n18596;
  assign n18598 =  a[17]  & ~n18597;
  assign n18599 = ~ a[17]  & n18597;
  assign n18600 = ~n18598 & ~n18599;
  assign n18601 = n18589 & ~n18600;
  assign n18602 = n18102 & n18274;
  assign n18603 = ~n18275 & ~n18602;
  assign n18604 = n6233 & n12537;
  assign n18605 = n5663 & n12543;
  assign n18606 = n5939 & n12540;
  assign n18607 = ~n18605 & ~n18606;
  assign n18608 = ~n18604 & n18607;
  assign n18609 = ~n5666 & n18608;
  assign n18610 = n15385 & n18608;
  assign n18611 = ~n18609 & ~n18610;
  assign n18612 =  a[17]  & ~n18611;
  assign n18613 = ~ a[17]  & n18611;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = n18603 & ~n18614;
  assign n18616 = n6233 & n12540;
  assign n18617 = n5663 & n12546;
  assign n18618 = n5939 & n12543;
  assign n18619 = ~n18617 & ~n18618;
  assign n18620 = ~n18616 & n18619;
  assign n18621 = n5666 & ~n15708;
  assign n18622 = n18620 & ~n18621;
  assign n18623 =  a[17]  & ~n18622;
  assign n18624 = ~n18622 & ~n18623;
  assign n18625 =  a[17]  & ~n18623;
  assign n18626 = ~n18624 & ~n18625;
  assign n18627 = n18270 & ~n18272;
  assign n18628 = ~n18273 & ~n18627;
  assign n18629 = ~n18626 & n18628;
  assign n18630 = ~n18626 & ~n18629;
  assign n18631 = n18628 & ~n18629;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = n6233 & n12543;
  assign n18634 = n5663 & n12549;
  assign n18635 = n5939 & n12546;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = ~n18633 & n18636;
  assign n18638 = n5666 & n15724;
  assign n18639 = n18637 & ~n18638;
  assign n18640 =  a[17]  & ~n18639;
  assign n18641 = ~n18639 & ~n18640;
  assign n18642 =  a[17]  & ~n18640;
  assign n18643 = ~n18641 & ~n18642;
  assign n18644 = ~n18265 & ~n18269;
  assign n18645 = ~n18268 & ~n18269;
  assign n18646 = ~n18644 & ~n18645;
  assign n18647 = ~n18643 & ~n18646;
  assign n18648 = ~n18643 & ~n18647;
  assign n18649 = ~n18646 & ~n18647;
  assign n18650 = ~n18648 & ~n18649;
  assign n18651 = n6233 & n12546;
  assign n18652 = n5663 & n12552;
  assign n18653 = n5939 & n12549;
  assign n18654 = ~n18652 & ~n18653;
  assign n18655 = ~n18651 & n18654;
  assign n18656 = n5666 & ~n15356;
  assign n18657 = n18655 & ~n18656;
  assign n18658 =  a[17]  & ~n18657;
  assign n18659 = ~n18657 & ~n18658;
  assign n18660 =  a[17]  & ~n18658;
  assign n18661 = ~n18659 & ~n18660;
  assign n18662 = ~n18260 & ~n18264;
  assign n18663 = ~n18263 & ~n18264;
  assign n18664 = ~n18662 & ~n18663;
  assign n18665 = ~n18661 & ~n18664;
  assign n18666 = ~n18661 & ~n18665;
  assign n18667 = ~n18664 & ~n18665;
  assign n18668 = ~n18666 & ~n18667;
  assign n18669 = n18161 & n18258;
  assign n18670 = ~n18259 & ~n18669;
  assign n18671 = n6233 & n12549;
  assign n18672 = n5663 & n12555;
  assign n18673 = n5939 & n12552;
  assign n18674 = ~n18672 & ~n18673;
  assign n18675 = ~n18671 & n18674;
  assign n18676 = ~n5666 & n18675;
  assign n18677 = ~n15764 & n18675;
  assign n18678 = ~n18676 & ~n18677;
  assign n18679 =  a[17]  & ~n18678;
  assign n18680 = ~ a[17]  & n18678;
  assign n18681 = ~n18679 & ~n18680;
  assign n18682 = n18670 & ~n18681;
  assign n18683 = n18254 & ~n18256;
  assign n18684 = ~n18257 & ~n18683;
  assign n18685 = n6233 & n12552;
  assign n18686 = n5663 & n12558;
  assign n18687 = n5939 & n12555;
  assign n18688 = ~n18686 & ~n18687;
  assign n18689 = ~n18685 & n18688;
  assign n18690 = ~n5666 & n18689;
  assign n18691 = n15791 & n18689;
  assign n18692 = ~n18690 & ~n18691;
  assign n18693 =  a[17]  & ~n18692;
  assign n18694 = ~ a[17]  & n18692;
  assign n18695 = ~n18693 & ~n18694;
  assign n18696 = n18684 & ~n18695;
  assign n18697 = n18193 & n18252;
  assign n18698 = ~n18253 & ~n18697;
  assign n18699 = n6233 & n12555;
  assign n18700 = n5663 & n12561;
  assign n18701 = n5939 & n12558;
  assign n18702 = ~n18700 & ~n18701;
  assign n18703 = ~n18699 & n18702;
  assign n18704 = ~n5666 & n18703;
  assign n18705 = n15816 & n18703;
  assign n18706 = ~n18704 & ~n18705;
  assign n18707 =  a[17]  & ~n18706;
  assign n18708 = ~ a[17]  & n18706;
  assign n18709 = ~n18707 & ~n18708;
  assign n18710 = n18698 & ~n18709;
  assign n18711 = n6233 & n12558;
  assign n18712 = n5663 & n12564;
  assign n18713 = n5939 & n12561;
  assign n18714 = ~n18712 & ~n18713;
  assign n18715 = ~n18711 & n18714;
  assign n18716 = n5666 & n15847;
  assign n18717 = n18715 & ~n18716;
  assign n18718 =  a[17]  & ~n18717;
  assign n18719 = ~n18717 & ~n18718;
  assign n18720 =  a[17]  & ~n18718;
  assign n18721 = ~n18719 & ~n18720;
  assign n18722 = n18248 & ~n18250;
  assign n18723 = ~n18251 & ~n18722;
  assign n18724 = ~n18721 & n18723;
  assign n18725 = ~n18721 & ~n18724;
  assign n18726 = n18723 & ~n18724;
  assign n18727 = ~n18725 & ~n18726;
  assign n18728 = ~n18235 & ~n18247;
  assign n18729 = ~n18246 & ~n18247;
  assign n18730 = ~n18728 & ~n18729;
  assign n18731 = n6233 & n12561;
  assign n18732 = n5663 & n12567;
  assign n18733 = n5939 & n12564;
  assign n18734 = ~n18732 & ~n18733;
  assign n18735 = ~n18731 & n18734;
  assign n18736 = ~n5666 & n18735;
  assign n18737 = n15905 & n18735;
  assign n18738 = ~n18736 & ~n18737;
  assign n18739 =  a[17]  & ~n18738;
  assign n18740 = ~ a[17]  & n18738;
  assign n18741 = ~n18739 & ~n18740;
  assign n18742 = ~n18730 & ~n18741;
  assign n18743 = n6233 & n12564;
  assign n18744 = n5663 & n12571;
  assign n18745 = n5939 & n12567;
  assign n18746 = ~n18744 & ~n18745;
  assign n18747 = ~n18743 & n18746;
  assign n18748 = n5666 & ~n15944;
  assign n18749 = n18747 & ~n18748;
  assign n18750 =  a[17]  & ~n18749;
  assign n18751 = ~n18749 & ~n18750;
  assign n18752 =  a[17]  & ~n18750;
  assign n18753 = ~n18751 & ~n18752;
  assign n18754 = ~n18219 & n18230;
  assign n18755 = ~n18231 & ~n18754;
  assign n18756 = ~n18753 & n18755;
  assign n18757 = ~n18753 & ~n18756;
  assign n18758 = n18755 & ~n18756;
  assign n18759 = ~n18757 & ~n18758;
  assign n18760 = n18216 & ~n18218;
  assign n18761 = ~n18219 & ~n18760;
  assign n18762 = n6233 & n12567;
  assign n18763 = n5663 & n12574;
  assign n18764 = n5939 & n12571;
  assign n18765 = ~n18763 & ~n18764;
  assign n18766 = ~n18762 & n18765;
  assign n18767 = ~n5666 & n18766;
  assign n18768 = ~n15989 & n18766;
  assign n18769 = ~n18767 & ~n18768;
  assign n18770 =  a[17]  & ~n18769;
  assign n18771 = ~ a[17]  & n18769;
  assign n18772 = ~n18770 & ~n18771;
  assign n18773 = n18761 & ~n18772;
  assign n18774 = n5939 & ~n12581;
  assign n18775 = n6233 & n12577;
  assign n18776 = ~n18774 & ~n18775;
  assign n18777 = n5666 & ~n16085;
  assign n18778 = n18776 & ~n18777;
  assign n18779 =  a[17]  & ~n18778;
  assign n18780 =  a[17]  & ~n18779;
  assign n18781 = ~n18778 & ~n18779;
  assign n18782 = ~n18780 & ~n18781;
  assign n18783 = ~n5658 & ~n12581;
  assign n18784 =  a[17]  & ~n18783;
  assign n18785 = ~n18782 & n18784;
  assign n18786 = n6233 & n12574;
  assign n18787 = n5663 & ~n12581;
  assign n18788 = n5939 & n12577;
  assign n18789 = ~n18787 & ~n18788;
  assign n18790 = ~n18786 & n18789;
  assign n18791 = ~n5666 & n18790;
  assign n18792 = n16094 & n18790;
  assign n18793 = ~n18791 & ~n18792;
  assign n18794 =  a[17]  & ~n18793;
  assign n18795 = ~ a[17]  & n18793;
  assign n18796 = ~n18794 & ~n18795;
  assign n18797 = n18785 & ~n18796;
  assign n18798 = n18217 & n18797;
  assign n18799 = n18797 & ~n18798;
  assign n18800 = n18217 & ~n18798;
  assign n18801 = ~n18799 & ~n18800;
  assign n18802 = n6233 & n12571;
  assign n18803 = n5663 & n12577;
  assign n18804 = n5939 & n12574;
  assign n18805 = ~n18803 & ~n18804;
  assign n18806 = ~n18802 & n18805;
  assign n18807 = n5666 & n16013;
  assign n18808 = n18806 & ~n18807;
  assign n18809 =  a[17]  & ~n18808;
  assign n18810 =  a[17]  & ~n18809;
  assign n18811 = ~n18808 & ~n18809;
  assign n18812 = ~n18810 & ~n18811;
  assign n18813 = ~n18801 & ~n18812;
  assign n18814 = ~n18798 & ~n18813;
  assign n18815 = ~n18761 & n18772;
  assign n18816 = ~n18773 & ~n18815;
  assign n18817 = ~n18814 & n18816;
  assign n18818 = ~n18773 & ~n18817;
  assign n18819 = ~n18759 & ~n18818;
  assign n18820 = ~n18756 & ~n18819;
  assign n18821 = n18730 & n18741;
  assign n18822 = ~n18742 & ~n18821;
  assign n18823 = ~n18820 & n18822;
  assign n18824 = ~n18742 & ~n18823;
  assign n18825 = ~n18727 & ~n18824;
  assign n18826 = ~n18724 & ~n18825;
  assign n18827 = n18698 & ~n18710;
  assign n18828 = ~n18709 & ~n18710;
  assign n18829 = ~n18827 & ~n18828;
  assign n18830 = ~n18826 & ~n18829;
  assign n18831 = ~n18710 & ~n18830;
  assign n18832 = n18684 & ~n18696;
  assign n18833 = ~n18695 & ~n18696;
  assign n18834 = ~n18832 & ~n18833;
  assign n18835 = ~n18831 & ~n18834;
  assign n18836 = ~n18696 & ~n18835;
  assign n18837 = ~n18670 & n18681;
  assign n18838 = ~n18682 & ~n18837;
  assign n18839 = ~n18836 & n18838;
  assign n18840 = ~n18682 & ~n18839;
  assign n18841 = ~n18668 & ~n18840;
  assign n18842 = ~n18665 & ~n18841;
  assign n18843 = ~n18650 & ~n18842;
  assign n18844 = ~n18647 & ~n18843;
  assign n18845 = ~n18632 & ~n18844;
  assign n18846 = ~n18629 & ~n18845;
  assign n18847 = n18603 & ~n18615;
  assign n18848 = ~n18614 & ~n18615;
  assign n18849 = ~n18847 & ~n18848;
  assign n18850 = ~n18846 & ~n18849;
  assign n18851 = ~n18615 & ~n18850;
  assign n18852 = ~n18589 & n18600;
  assign n18853 = ~n18601 & ~n18852;
  assign n18854 = ~n18851 & n18853;
  assign n18855 = ~n18601 & ~n18854;
  assign n18856 = ~n18587 & ~n18855;
  assign n18857 = ~n18584 & ~n18856;
  assign n18858 = ~n18569 & ~n18857;
  assign n18859 = ~n18566 & ~n18858;
  assign n18860 = ~n18551 & ~n18859;
  assign n18861 = ~n18548 & ~n18860;
  assign n18862 = ~n18533 & ~n18861;
  assign n18863 = ~n18530 & ~n18862;
  assign n18864 = ~n18515 & ~n18863;
  assign n18865 = ~n18512 & ~n18864;
  assign n18866 = ~n18497 & ~n18865;
  assign n18867 = ~n18494 & ~n18866;
  assign n18868 = ~n18479 & ~n18867;
  assign n18869 = ~n18476 & ~n18868;
  assign n18870 = ~n18461 & ~n18869;
  assign n18871 = ~n18458 & ~n18870;
  assign n18872 = ~n18443 & ~n18871;
  assign n18873 = ~n18440 & ~n18872;
  assign n18874 = ~n18425 & ~n18873;
  assign n18875 = ~n18422 & ~n18874;
  assign n18876 = ~n18408 & ~n18875;
  assign n18877 = n18408 & n18875;
  assign n18878 = ~n18876 & ~n18877;
  assign n18879 = n7101 & n12889;
  assign n18880 = n6402 & n12502;
  assign n18881 = n6951 & n12769;
  assign n18882 = ~n18880 & ~n18881;
  assign n18883 = ~n18879 & n18882;
  assign n18884 = n6397 & n12895;
  assign n18885 = n18883 & ~n18884;
  assign n18886 =  a[14]  & ~n18885;
  assign n18887 =  a[14]  & ~n18886;
  assign n18888 = ~n18885 & ~n18886;
  assign n18889 = ~n18887 & ~n18888;
  assign n18890 = n18878 & ~n18889;
  assign n18891 = ~n18876 & ~n18890;
  assign n18892 = ~n18405 & ~n18891;
  assign n18893 = n18405 & n18891;
  assign n18894 = ~n18892 & ~n18893;
  assign n18895 = n7983 & n13515;
  assign n18896 = n7291 & n13518;
  assign n18897 = n7632 & n13521;
  assign n18898 = ~n18896 & ~n18897;
  assign n18899 = ~n18895 & n18898;
  assign n18900 = n7294 & n13541;
  assign n18901 = n18899 & ~n18900;
  assign n18902 =  a[11]  & ~n18901;
  assign n18903 =  a[11]  & ~n18902;
  assign n18904 = ~n18901 & ~n18902;
  assign n18905 = ~n18903 & ~n18904;
  assign n18906 = n18894 & ~n18905;
  assign n18907 = ~n18892 & ~n18906;
  assign n18908 = ~n18402 & ~n18907;
  assign n18909 = n18402 & n18907;
  assign n18910 = ~n18908 & ~n18909;
  assign n18911 = n9331 & ~n13627;
  assign n18912 = n8418 & n13630;
  assign n18913 = n8860 & n13633;
  assign n18914 = ~n18912 & ~n18913;
  assign n18915 = ~n18911 & n18914;
  assign n18916 = n8421 & ~n13654;
  assign n18917 = n18915 & ~n18916;
  assign n18918 =  a[8]  & ~n18917;
  assign n18919 =  a[8]  & ~n18918;
  assign n18920 = ~n18917 & ~n18918;
  assign n18921 = ~n18919 & ~n18920;
  assign n18922 = n18910 & ~n18921;
  assign n18923 = ~n18908 & ~n18922;
  assign n18924 = n9331 & n13941;
  assign n18925 = n8418 & n13633;
  assign n18926 = n8860 & ~n13627;
  assign n18927 = ~n18925 & ~n18926;
  assign n18928 = ~n18924 & n18927;
  assign n18929 = n8421 & n14136;
  assign n18930 = n18928 & ~n18929;
  assign n18931 =  a[8]  & ~n18930;
  assign n18932 =  a[8]  & ~n18931;
  assign n18933 = ~n18930 & ~n18931;
  assign n18934 = ~n18932 & ~n18933;
  assign n18935 = ~n18923 & ~n18934;
  assign n18936 = ~n18923 & ~n18935;
  assign n18937 = ~n18934 & ~n18935;
  assign n18938 = ~n18936 & ~n18937;
  assign n18939 = n17918 & n18375;
  assign n18940 = ~n18376 & ~n18939;
  assign n18941 = ~n18938 & n18940;
  assign n18942 = ~n18935 & ~n18941;
  assign n18943 = ~n18399 & ~n18942;
  assign n18944 = ~n18399 & ~n18943;
  assign n18945 = ~n18942 & ~n18943;
  assign n18946 = ~n18944 & ~n18945;
  assign n18947 = n18894 & ~n18906;
  assign n18948 = ~n18905 & ~n18906;
  assign n18949 = ~n18947 & ~n18948;
  assign n18950 = n18878 & ~n18890;
  assign n18951 = ~n18889 & ~n18890;
  assign n18952 = ~n18950 & ~n18951;
  assign n18953 = n18425 & n18873;
  assign n18954 = ~n18874 & ~n18953;
  assign n18955 = n7101 & n12769;
  assign n18956 = n6402 & n12370;
  assign n18957 = n6951 & n12502;
  assign n18958 = ~n18956 & ~n18957;
  assign n18959 = ~n18955 & n18958;
  assign n18960 = ~n6397 & n18959;
  assign n18961 = ~n12999 & n18959;
  assign n18962 = ~n18960 & ~n18961;
  assign n18963 =  a[14]  & ~n18962;
  assign n18964 = ~ a[14]  & n18962;
  assign n18965 = ~n18963 & ~n18964;
  assign n18966 = n18954 & ~n18965;
  assign n18967 = n18443 & n18871;
  assign n18968 = ~n18872 & ~n18967;
  assign n18969 = n7101 & n12502;
  assign n18970 = n6402 & n12505;
  assign n18971 = n6951 & n12370;
  assign n18972 = ~n18970 & ~n18971;
  assign n18973 = ~n18969 & n18972;
  assign n18974 = ~n6397 & n18973;
  assign n18975 = n13736 & n18973;
  assign n18976 = ~n18974 & ~n18975;
  assign n18977 =  a[14]  & ~n18976;
  assign n18978 = ~ a[14]  & n18976;
  assign n18979 = ~n18977 & ~n18978;
  assign n18980 = n18968 & ~n18979;
  assign n18981 = n18461 & n18869;
  assign n18982 = ~n18870 & ~n18981;
  assign n18983 = n7101 & n12370;
  assign n18984 = n6402 & n12508;
  assign n18985 = n6951 & n12505;
  assign n18986 = ~n18984 & ~n18985;
  assign n18987 = ~n18983 & n18986;
  assign n18988 = ~n6397 & n18987;
  assign n18989 = n13748 & n18987;
  assign n18990 = ~n18988 & ~n18989;
  assign n18991 =  a[14]  & ~n18990;
  assign n18992 = ~ a[14]  & n18990;
  assign n18993 = ~n18991 & ~n18992;
  assign n18994 = n18982 & ~n18993;
  assign n18995 = n18479 & n18867;
  assign n18996 = ~n18868 & ~n18995;
  assign n18997 = n7101 & n12505;
  assign n18998 = n6402 & n12513;
  assign n18999 = n6951 & n12508;
  assign n19000 = ~n18998 & ~n18999;
  assign n19001 = ~n18997 & n19000;
  assign n19002 = ~n6397 & n19001;
  assign n19003 = n14051 & n19001;
  assign n19004 = ~n19002 & ~n19003;
  assign n19005 =  a[14]  & ~n19004;
  assign n19006 = ~ a[14]  & n19004;
  assign n19007 = ~n19005 & ~n19006;
  assign n19008 = n18996 & ~n19007;
  assign n19009 = n18497 & n18865;
  assign n19010 = ~n18866 & ~n19009;
  assign n19011 = n7101 & n12508;
  assign n19012 = n6402 & n12511;
  assign n19013 = n6951 & n12513;
  assign n19014 = ~n19012 & ~n19013;
  assign n19015 = ~n19011 & n19014;
  assign n19016 = ~n6397 & n19015;
  assign n19017 = ~n13863 & n19015;
  assign n19018 = ~n19016 & ~n19017;
  assign n19019 =  a[14]  & ~n19018;
  assign n19020 = ~ a[14]  & n19018;
  assign n19021 = ~n19019 & ~n19020;
  assign n19022 = n19010 & ~n19021;
  assign n19023 = n18515 & n18863;
  assign n19024 = ~n18864 & ~n19023;
  assign n19025 = n7101 & n12513;
  assign n19026 = n6402 & n12516;
  assign n19027 = n6951 & n12511;
  assign n19028 = ~n19026 & ~n19027;
  assign n19029 = ~n19025 & n19028;
  assign n19030 = ~n6397 & n19029;
  assign n19031 = ~n14177 & n19029;
  assign n19032 = ~n19030 & ~n19031;
  assign n19033 =  a[14]  & ~n19032;
  assign n19034 = ~ a[14]  & n19032;
  assign n19035 = ~n19033 & ~n19034;
  assign n19036 = n19024 & ~n19035;
  assign n19037 = n18533 & n18861;
  assign n19038 = ~n18862 & ~n19037;
  assign n19039 = n7101 & n12511;
  assign n19040 = n6402 & n12519;
  assign n19041 = n6951 & n12516;
  assign n19042 = ~n19040 & ~n19041;
  assign n19043 = ~n19039 & n19042;
  assign n19044 = ~n6397 & n19043;
  assign n19045 = n14233 & n19043;
  assign n19046 = ~n19044 & ~n19045;
  assign n19047 =  a[14]  & ~n19046;
  assign n19048 = ~ a[14]  & n19046;
  assign n19049 = ~n19047 & ~n19048;
  assign n19050 = n19038 & ~n19049;
  assign n19051 = n18551 & n18859;
  assign n19052 = ~n18860 & ~n19051;
  assign n19053 = n7101 & n12516;
  assign n19054 = n6402 & n12522;
  assign n19055 = n6951 & n12519;
  assign n19056 = ~n19054 & ~n19055;
  assign n19057 = ~n19053 & n19056;
  assign n19058 = ~n6397 & n19057;
  assign n19059 = n14443 & n19057;
  assign n19060 = ~n19058 & ~n19059;
  assign n19061 =  a[14]  & ~n19060;
  assign n19062 = ~ a[14]  & n19060;
  assign n19063 = ~n19061 & ~n19062;
  assign n19064 = n19052 & ~n19063;
  assign n19065 = n18569 & n18857;
  assign n19066 = ~n18858 & ~n19065;
  assign n19067 = n7101 & n12519;
  assign n19068 = n6402 & n12525;
  assign n19069 = n6951 & n12522;
  assign n19070 = ~n19068 & ~n19069;
  assign n19071 = ~n19067 & n19070;
  assign n19072 = ~n6397 & n19071;
  assign n19073 = ~n14454 & n19071;
  assign n19074 = ~n19072 & ~n19073;
  assign n19075 =  a[14]  & ~n19074;
  assign n19076 = ~ a[14]  & n19074;
  assign n19077 = ~n19075 & ~n19076;
  assign n19078 = n19066 & ~n19077;
  assign n19079 = n18587 & n18855;
  assign n19080 = ~n18856 & ~n19079;
  assign n19081 = n7101 & n12522;
  assign n19082 = n6402 & n12528;
  assign n19083 = n6951 & n12525;
  assign n19084 = ~n19082 & ~n19083;
  assign n19085 = ~n19081 & n19084;
  assign n19086 = ~n6397 & n19085;
  assign n19087 = ~n14837 & n19085;
  assign n19088 = ~n19086 & ~n19087;
  assign n19089 =  a[14]  & ~n19088;
  assign n19090 = ~ a[14]  & n19088;
  assign n19091 = ~n19089 & ~n19090;
  assign n19092 = n19080 & ~n19091;
  assign n19093 = n7101 & n12525;
  assign n19094 = n6402 & n12531;
  assign n19095 = n6951 & n12528;
  assign n19096 = ~n19094 & ~n19095;
  assign n19097 = ~n19093 & n19096;
  assign n19098 = n6397 & n14608;
  assign n19099 = n19097 & ~n19098;
  assign n19100 =  a[14]  & ~n19099;
  assign n19101 = ~n19099 & ~n19100;
  assign n19102 =  a[14]  & ~n19100;
  assign n19103 = ~n19101 & ~n19102;
  assign n19104 = n18851 & ~n18853;
  assign n19105 = ~n18854 & ~n19104;
  assign n19106 = ~n19103 & n19105;
  assign n19107 = ~n19103 & ~n19106;
  assign n19108 = n19105 & ~n19106;
  assign n19109 = ~n19107 & ~n19108;
  assign n19110 = n7101 & n12528;
  assign n19111 = n6402 & n12534;
  assign n19112 = n6951 & n12531;
  assign n19113 = ~n19111 & ~n19112;
  assign n19114 = ~n19110 & n19113;
  assign n19115 = n6397 & ~n15003;
  assign n19116 = n19114 & ~n19115;
  assign n19117 =  a[14]  & ~n19116;
  assign n19118 = ~n19116 & ~n19117;
  assign n19119 =  a[14]  & ~n19117;
  assign n19120 = ~n19118 & ~n19119;
  assign n19121 = ~n18846 & ~n18850;
  assign n19122 = ~n18849 & ~n18850;
  assign n19123 = ~n19121 & ~n19122;
  assign n19124 = ~n19120 & ~n19123;
  assign n19125 = ~n19120 & ~n19124;
  assign n19126 = ~n19123 & ~n19124;
  assign n19127 = ~n19125 & ~n19126;
  assign n19128 = n18632 & n18844;
  assign n19129 = ~n18845 & ~n19128;
  assign n19130 = n7101 & n12531;
  assign n19131 = n6402 & n12537;
  assign n19132 = n6951 & n12534;
  assign n19133 = ~n19131 & ~n19132;
  assign n19134 = ~n19130 & n19133;
  assign n19135 = ~n6397 & n19134;
  assign n19136 = ~n15255 & n19134;
  assign n19137 = ~n19135 & ~n19136;
  assign n19138 =  a[14]  & ~n19137;
  assign n19139 = ~ a[14]  & n19137;
  assign n19140 = ~n19138 & ~n19139;
  assign n19141 = n19129 & ~n19140;
  assign n19142 = n18650 & n18842;
  assign n19143 = ~n18843 & ~n19142;
  assign n19144 = n7101 & n12534;
  assign n19145 = n6402 & n12540;
  assign n19146 = n6951 & n12537;
  assign n19147 = ~n19145 & ~n19146;
  assign n19148 = ~n19144 & n19147;
  assign n19149 = ~n6397 & n19148;
  assign n19150 = n15096 & n19148;
  assign n19151 = ~n19149 & ~n19150;
  assign n19152 =  a[14]  & ~n19151;
  assign n19153 = ~ a[14]  & n19151;
  assign n19154 = ~n19152 & ~n19153;
  assign n19155 = n19143 & ~n19154;
  assign n19156 = n18668 & n18840;
  assign n19157 = ~n18841 & ~n19156;
  assign n19158 = n7101 & n12537;
  assign n19159 = n6402 & n12543;
  assign n19160 = n6951 & n12540;
  assign n19161 = ~n19159 & ~n19160;
  assign n19162 = ~n19158 & n19161;
  assign n19163 = ~n6397 & n19162;
  assign n19164 = n15385 & n19162;
  assign n19165 = ~n19163 & ~n19164;
  assign n19166 =  a[14]  & ~n19165;
  assign n19167 = ~ a[14]  & n19165;
  assign n19168 = ~n19166 & ~n19167;
  assign n19169 = n19157 & ~n19168;
  assign n19170 = n7101 & n12540;
  assign n19171 = n6402 & n12546;
  assign n19172 = n6951 & n12543;
  assign n19173 = ~n19171 & ~n19172;
  assign n19174 = ~n19170 & n19173;
  assign n19175 = n6397 & ~n15708;
  assign n19176 = n19174 & ~n19175;
  assign n19177 =  a[14]  & ~n19176;
  assign n19178 = ~n19176 & ~n19177;
  assign n19179 =  a[14]  & ~n19177;
  assign n19180 = ~n19178 & ~n19179;
  assign n19181 = n18836 & ~n18838;
  assign n19182 = ~n18839 & ~n19181;
  assign n19183 = ~n19180 & n19182;
  assign n19184 = ~n19180 & ~n19183;
  assign n19185 = n19182 & ~n19183;
  assign n19186 = ~n19184 & ~n19185;
  assign n19187 = n7101 & n12543;
  assign n19188 = n6402 & n12549;
  assign n19189 = n6951 & n12546;
  assign n19190 = ~n19188 & ~n19189;
  assign n19191 = ~n19187 & n19190;
  assign n19192 = n6397 & n15724;
  assign n19193 = n19191 & ~n19192;
  assign n19194 =  a[14]  & ~n19193;
  assign n19195 = ~n19193 & ~n19194;
  assign n19196 =  a[14]  & ~n19194;
  assign n19197 = ~n19195 & ~n19196;
  assign n19198 = ~n18831 & ~n18835;
  assign n19199 = ~n18834 & ~n18835;
  assign n19200 = ~n19198 & ~n19199;
  assign n19201 = ~n19197 & ~n19200;
  assign n19202 = ~n19197 & ~n19201;
  assign n19203 = ~n19200 & ~n19201;
  assign n19204 = ~n19202 & ~n19203;
  assign n19205 = n7101 & n12546;
  assign n19206 = n6402 & n12552;
  assign n19207 = n6951 & n12549;
  assign n19208 = ~n19206 & ~n19207;
  assign n19209 = ~n19205 & n19208;
  assign n19210 = n6397 & ~n15356;
  assign n19211 = n19209 & ~n19210;
  assign n19212 =  a[14]  & ~n19211;
  assign n19213 = ~n19211 & ~n19212;
  assign n19214 =  a[14]  & ~n19212;
  assign n19215 = ~n19213 & ~n19214;
  assign n19216 = ~n18826 & ~n18830;
  assign n19217 = ~n18829 & ~n18830;
  assign n19218 = ~n19216 & ~n19217;
  assign n19219 = ~n19215 & ~n19218;
  assign n19220 = ~n19215 & ~n19219;
  assign n19221 = ~n19218 & ~n19219;
  assign n19222 = ~n19220 & ~n19221;
  assign n19223 = n18727 & n18824;
  assign n19224 = ~n18825 & ~n19223;
  assign n19225 = n7101 & n12549;
  assign n19226 = n6402 & n12555;
  assign n19227 = n6951 & n12552;
  assign n19228 = ~n19226 & ~n19227;
  assign n19229 = ~n19225 & n19228;
  assign n19230 = ~n6397 & n19229;
  assign n19231 = ~n15764 & n19229;
  assign n19232 = ~n19230 & ~n19231;
  assign n19233 =  a[14]  & ~n19232;
  assign n19234 = ~ a[14]  & n19232;
  assign n19235 = ~n19233 & ~n19234;
  assign n19236 = n19224 & ~n19235;
  assign n19237 = n18820 & ~n18822;
  assign n19238 = ~n18823 & ~n19237;
  assign n19239 = n7101 & n12552;
  assign n19240 = n6402 & n12558;
  assign n19241 = n6951 & n12555;
  assign n19242 = ~n19240 & ~n19241;
  assign n19243 = ~n19239 & n19242;
  assign n19244 = ~n6397 & n19243;
  assign n19245 = n15791 & n19243;
  assign n19246 = ~n19244 & ~n19245;
  assign n19247 =  a[14]  & ~n19246;
  assign n19248 = ~ a[14]  & n19246;
  assign n19249 = ~n19247 & ~n19248;
  assign n19250 = n19238 & ~n19249;
  assign n19251 = n18759 & n18818;
  assign n19252 = ~n18819 & ~n19251;
  assign n19253 = n7101 & n12555;
  assign n19254 = n6402 & n12561;
  assign n19255 = n6951 & n12558;
  assign n19256 = ~n19254 & ~n19255;
  assign n19257 = ~n19253 & n19256;
  assign n19258 = ~n6397 & n19257;
  assign n19259 = n15816 & n19257;
  assign n19260 = ~n19258 & ~n19259;
  assign n19261 =  a[14]  & ~n19260;
  assign n19262 = ~ a[14]  & n19260;
  assign n19263 = ~n19261 & ~n19262;
  assign n19264 = n19252 & ~n19263;
  assign n19265 = n7101 & n12558;
  assign n19266 = n6402 & n12564;
  assign n19267 = n6951 & n12561;
  assign n19268 = ~n19266 & ~n19267;
  assign n19269 = ~n19265 & n19268;
  assign n19270 = n6397 & n15847;
  assign n19271 = n19269 & ~n19270;
  assign n19272 =  a[14]  & ~n19271;
  assign n19273 = ~n19271 & ~n19272;
  assign n19274 =  a[14]  & ~n19272;
  assign n19275 = ~n19273 & ~n19274;
  assign n19276 = n18814 & ~n18816;
  assign n19277 = ~n18817 & ~n19276;
  assign n19278 = ~n19275 & n19277;
  assign n19279 = ~n19275 & ~n19278;
  assign n19280 = n19277 & ~n19278;
  assign n19281 = ~n19279 & ~n19280;
  assign n19282 = ~n18801 & ~n18813;
  assign n19283 = ~n18812 & ~n18813;
  assign n19284 = ~n19282 & ~n19283;
  assign n19285 = n7101 & n12561;
  assign n19286 = n6402 & n12567;
  assign n19287 = n6951 & n12564;
  assign n19288 = ~n19286 & ~n19287;
  assign n19289 = ~n19285 & n19288;
  assign n19290 = ~n6397 & n19289;
  assign n19291 = n15905 & n19289;
  assign n19292 = ~n19290 & ~n19291;
  assign n19293 =  a[14]  & ~n19292;
  assign n19294 = ~ a[14]  & n19292;
  assign n19295 = ~n19293 & ~n19294;
  assign n19296 = ~n19284 & ~n19295;
  assign n19297 = n7101 & n12564;
  assign n19298 = n6402 & n12571;
  assign n19299 = n6951 & n12567;
  assign n19300 = ~n19298 & ~n19299;
  assign n19301 = ~n19297 & n19300;
  assign n19302 = n6397 & ~n15944;
  assign n19303 = n19301 & ~n19302;
  assign n19304 =  a[14]  & ~n19303;
  assign n19305 = ~n19303 & ~n19304;
  assign n19306 =  a[14]  & ~n19304;
  assign n19307 = ~n19305 & ~n19306;
  assign n19308 = ~n18785 & n18796;
  assign n19309 = ~n18797 & ~n19308;
  assign n19310 = ~n19307 & n19309;
  assign n19311 = ~n19307 & ~n19310;
  assign n19312 = n19309 & ~n19310;
  assign n19313 = ~n19311 & ~n19312;
  assign n19314 = n18782 & ~n18784;
  assign n19315 = ~n18785 & ~n19314;
  assign n19316 = n7101 & n12567;
  assign n19317 = n6402 & n12574;
  assign n19318 = n6951 & n12571;
  assign n19319 = ~n19317 & ~n19318;
  assign n19320 = ~n19316 & n19319;
  assign n19321 = ~n6397 & n19320;
  assign n19322 = ~n15989 & n19320;
  assign n19323 = ~n19321 & ~n19322;
  assign n19324 =  a[14]  & ~n19323;
  assign n19325 = ~ a[14]  & n19323;
  assign n19326 = ~n19324 & ~n19325;
  assign n19327 = n19315 & ~n19326;
  assign n19328 = n6951 & ~n12581;
  assign n19329 = n7101 & n12577;
  assign n19330 = ~n19328 & ~n19329;
  assign n19331 = n6397 & ~n16085;
  assign n19332 = n19330 & ~n19331;
  assign n19333 =  a[14]  & ~n19332;
  assign n19334 =  a[14]  & ~n19333;
  assign n19335 = ~n19332 & ~n19333;
  assign n19336 = ~n19334 & ~n19335;
  assign n19337 = ~n6393 & ~n12581;
  assign n19338 =  a[14]  & ~n19337;
  assign n19339 = ~n19336 & n19338;
  assign n19340 = n7101 & n12574;
  assign n19341 = n6402 & ~n12581;
  assign n19342 = n6951 & n12577;
  assign n19343 = ~n19341 & ~n19342;
  assign n19344 = ~n19340 & n19343;
  assign n19345 = ~n6397 & n19344;
  assign n19346 = n16094 & n19344;
  assign n19347 = ~n19345 & ~n19346;
  assign n19348 =  a[14]  & ~n19347;
  assign n19349 = ~ a[14]  & n19347;
  assign n19350 = ~n19348 & ~n19349;
  assign n19351 = n19339 & ~n19350;
  assign n19352 = n18783 & n19351;
  assign n19353 = n19351 & ~n19352;
  assign n19354 = n18783 & ~n19352;
  assign n19355 = ~n19353 & ~n19354;
  assign n19356 = n7101 & n12571;
  assign n19357 = n6402 & n12577;
  assign n19358 = n6951 & n12574;
  assign n19359 = ~n19357 & ~n19358;
  assign n19360 = ~n19356 & n19359;
  assign n19361 = n6397 & n16013;
  assign n19362 = n19360 & ~n19361;
  assign n19363 =  a[14]  & ~n19362;
  assign n19364 =  a[14]  & ~n19363;
  assign n19365 = ~n19362 & ~n19363;
  assign n19366 = ~n19364 & ~n19365;
  assign n19367 = ~n19355 & ~n19366;
  assign n19368 = ~n19352 & ~n19367;
  assign n19369 = ~n19315 & n19326;
  assign n19370 = ~n19327 & ~n19369;
  assign n19371 = ~n19368 & n19370;
  assign n19372 = ~n19327 & ~n19371;
  assign n19373 = ~n19313 & ~n19372;
  assign n19374 = ~n19310 & ~n19373;
  assign n19375 = n19284 & n19295;
  assign n19376 = ~n19296 & ~n19375;
  assign n19377 = ~n19374 & n19376;
  assign n19378 = ~n19296 & ~n19377;
  assign n19379 = ~n19281 & ~n19378;
  assign n19380 = ~n19278 & ~n19379;
  assign n19381 = n19252 & ~n19264;
  assign n19382 = ~n19263 & ~n19264;
  assign n19383 = ~n19381 & ~n19382;
  assign n19384 = ~n19380 & ~n19383;
  assign n19385 = ~n19264 & ~n19384;
  assign n19386 = n19238 & ~n19250;
  assign n19387 = ~n19249 & ~n19250;
  assign n19388 = ~n19386 & ~n19387;
  assign n19389 = ~n19385 & ~n19388;
  assign n19390 = ~n19250 & ~n19389;
  assign n19391 = ~n19224 & n19235;
  assign n19392 = ~n19236 & ~n19391;
  assign n19393 = ~n19390 & n19392;
  assign n19394 = ~n19236 & ~n19393;
  assign n19395 = ~n19222 & ~n19394;
  assign n19396 = ~n19219 & ~n19395;
  assign n19397 = ~n19204 & ~n19396;
  assign n19398 = ~n19201 & ~n19397;
  assign n19399 = ~n19186 & ~n19398;
  assign n19400 = ~n19183 & ~n19399;
  assign n19401 = n19157 & ~n19169;
  assign n19402 = ~n19168 & ~n19169;
  assign n19403 = ~n19401 & ~n19402;
  assign n19404 = ~n19400 & ~n19403;
  assign n19405 = ~n19169 & ~n19404;
  assign n19406 = n19143 & ~n19155;
  assign n19407 = ~n19154 & ~n19155;
  assign n19408 = ~n19406 & ~n19407;
  assign n19409 = ~n19405 & ~n19408;
  assign n19410 = ~n19155 & ~n19409;
  assign n19411 = ~n19129 & n19140;
  assign n19412 = ~n19141 & ~n19411;
  assign n19413 = ~n19410 & n19412;
  assign n19414 = ~n19141 & ~n19413;
  assign n19415 = ~n19127 & ~n19414;
  assign n19416 = ~n19124 & ~n19415;
  assign n19417 = ~n19109 & ~n19416;
  assign n19418 = ~n19106 & ~n19417;
  assign n19419 = n19080 & ~n19092;
  assign n19420 = ~n19091 & ~n19092;
  assign n19421 = ~n19419 & ~n19420;
  assign n19422 = ~n19418 & ~n19421;
  assign n19423 = ~n19092 & ~n19422;
  assign n19424 = n19066 & ~n19078;
  assign n19425 = ~n19077 & ~n19078;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = ~n19423 & ~n19426;
  assign n19428 = ~n19078 & ~n19427;
  assign n19429 = n19052 & ~n19064;
  assign n19430 = ~n19063 & ~n19064;
  assign n19431 = ~n19429 & ~n19430;
  assign n19432 = ~n19428 & ~n19431;
  assign n19433 = ~n19064 & ~n19432;
  assign n19434 = n19038 & ~n19050;
  assign n19435 = ~n19049 & ~n19050;
  assign n19436 = ~n19434 & ~n19435;
  assign n19437 = ~n19433 & ~n19436;
  assign n19438 = ~n19050 & ~n19437;
  assign n19439 = n19024 & ~n19036;
  assign n19440 = ~n19035 & ~n19036;
  assign n19441 = ~n19439 & ~n19440;
  assign n19442 = ~n19438 & ~n19441;
  assign n19443 = ~n19036 & ~n19442;
  assign n19444 = n19010 & ~n19022;
  assign n19445 = ~n19021 & ~n19022;
  assign n19446 = ~n19444 & ~n19445;
  assign n19447 = ~n19443 & ~n19446;
  assign n19448 = ~n19022 & ~n19447;
  assign n19449 = n18996 & ~n19008;
  assign n19450 = ~n19007 & ~n19008;
  assign n19451 = ~n19449 & ~n19450;
  assign n19452 = ~n19448 & ~n19451;
  assign n19453 = ~n19008 & ~n19452;
  assign n19454 = n18982 & ~n18994;
  assign n19455 = ~n18993 & ~n18994;
  assign n19456 = ~n19454 & ~n19455;
  assign n19457 = ~n19453 & ~n19456;
  assign n19458 = ~n18994 & ~n19457;
  assign n19459 = n18968 & ~n18980;
  assign n19460 = ~n18979 & ~n18980;
  assign n19461 = ~n19459 & ~n19460;
  assign n19462 = ~n19458 & ~n19461;
  assign n19463 = ~n18980 & ~n19462;
  assign n19464 = ~n18954 & n18965;
  assign n19465 = ~n18966 & ~n19464;
  assign n19466 = ~n19463 & n19465;
  assign n19467 = ~n18966 & ~n19466;
  assign n19468 = ~n18952 & ~n19467;
  assign n19469 = n18952 & n19467;
  assign n19470 = ~n19468 & ~n19469;
  assign n19471 = n7983 & n13521;
  assign n19472 = n7291 & n13491;
  assign n19473 = n7632 & n13518;
  assign n19474 = ~n19472 & ~n19473;
  assign n19475 = ~n19471 & n19474;
  assign n19476 = n7294 & ~n13909;
  assign n19477 = n19475 & ~n19476;
  assign n19478 =  a[11]  & ~n19477;
  assign n19479 =  a[11]  & ~n19478;
  assign n19480 = ~n19477 & ~n19478;
  assign n19481 = ~n19479 & ~n19480;
  assign n19482 = n19470 & ~n19481;
  assign n19483 = ~n19468 & ~n19482;
  assign n19484 = ~n18949 & ~n19483;
  assign n19485 = n18949 & n19483;
  assign n19486 = ~n19484 & ~n19485;
  assign n19487 = n9331 & n13633;
  assign n19488 = n8418 & n13597;
  assign n19489 = n8860 & n13630;
  assign n19490 = ~n19488 & ~n19489;
  assign n19491 = ~n19487 & n19490;
  assign n19492 = n8421 & n13929;
  assign n19493 = n19491 & ~n19492;
  assign n19494 =  a[8]  & ~n19493;
  assign n19495 =  a[8]  & ~n19494;
  assign n19496 = ~n19493 & ~n19494;
  assign n19497 = ~n19495 & ~n19496;
  assign n19498 = n19486 & ~n19497;
  assign n19499 = ~n19484 & ~n19498;
  assign n19500 = ~n13438 & ~n15076;
  assign n19501 = n9867 & n13941;
  assign n19502 = ~n19500 & ~n19501;
  assign n19503 = ~n9870 & n19502;
  assign n19504 = n13951 & n19502;
  assign n19505 = ~n19503 & ~n19504;
  assign n19506 =  a[5]  & ~n19505;
  assign n19507 = ~ a[5]  & n19505;
  assign n19508 = ~n19506 & ~n19507;
  assign n19509 = ~n19499 & ~n19508;
  assign n19510 = n18910 & ~n18922;
  assign n19511 = ~n18921 & ~n18922;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = n19499 & n19508;
  assign n19514 = ~n19509 & ~n19513;
  assign n19515 = ~n19512 & n19514;
  assign n19516 = ~n19509 & ~n19515;
  assign n19517 = n18938 & ~n18940;
  assign n19518 = ~n18941 & ~n19517;
  assign n19519 = ~n19516 & n19518;
  assign n19520 = ~n19512 & ~n19515;
  assign n19521 = n19514 & ~n19515;
  assign n19522 = ~n19520 & ~n19521;
  assign n19523 = n19486 & ~n19498;
  assign n19524 = ~n19497 & ~n19498;
  assign n19525 = ~n19523 & ~n19524;
  assign n19526 = n19470 & ~n19482;
  assign n19527 = ~n19481 & ~n19482;
  assign n19528 = ~n19526 & ~n19527;
  assign n19529 = n7983 & n13518;
  assign n19530 = n7291 & n12889;
  assign n19531 = n7632 & n13491;
  assign n19532 = ~n19530 & ~n19531;
  assign n19533 = ~n19529 & n19532;
  assign n19534 = n7294 & n13584;
  assign n19535 = n19533 & ~n19534;
  assign n19536 =  a[11]  & ~n19535;
  assign n19537 = ~n19535 & ~n19536;
  assign n19538 =  a[11]  & ~n19536;
  assign n19539 = ~n19537 & ~n19538;
  assign n19540 = n19463 & ~n19465;
  assign n19541 = ~n19466 & ~n19540;
  assign n19542 = ~n19539 & n19541;
  assign n19543 = ~n19539 & ~n19542;
  assign n19544 = n19541 & ~n19542;
  assign n19545 = ~n19543 & ~n19544;
  assign n19546 = n7983 & n13491;
  assign n19547 = n7291 & n12769;
  assign n19548 = n7632 & n12889;
  assign n19549 = ~n19547 & ~n19548;
  assign n19550 = ~n19546 & n19549;
  assign n19551 = n7294 & ~n13503;
  assign n19552 = n19550 & ~n19551;
  assign n19553 =  a[11]  & ~n19552;
  assign n19554 = ~n19552 & ~n19553;
  assign n19555 =  a[11]  & ~n19553;
  assign n19556 = ~n19554 & ~n19555;
  assign n19557 = ~n19458 & ~n19462;
  assign n19558 = ~n19461 & ~n19462;
  assign n19559 = ~n19557 & ~n19558;
  assign n19560 = ~n19556 & ~n19559;
  assign n19561 = ~n19556 & ~n19560;
  assign n19562 = ~n19559 & ~n19560;
  assign n19563 = ~n19561 & ~n19562;
  assign n19564 = n7983 & n12889;
  assign n19565 = n7291 & n12502;
  assign n19566 = n7632 & n12769;
  assign n19567 = ~n19565 & ~n19566;
  assign n19568 = ~n19564 & n19567;
  assign n19569 = n7294 & n12895;
  assign n19570 = n19568 & ~n19569;
  assign n19571 =  a[11]  & ~n19570;
  assign n19572 = ~n19570 & ~n19571;
  assign n19573 =  a[11]  & ~n19571;
  assign n19574 = ~n19572 & ~n19573;
  assign n19575 = ~n19453 & ~n19457;
  assign n19576 = ~n19456 & ~n19457;
  assign n19577 = ~n19575 & ~n19576;
  assign n19578 = ~n19574 & ~n19577;
  assign n19579 = ~n19574 & ~n19578;
  assign n19580 = ~n19577 & ~n19578;
  assign n19581 = ~n19579 & ~n19580;
  assign n19582 = n7983 & n12769;
  assign n19583 = n7291 & n12370;
  assign n19584 = n7632 & n12502;
  assign n19585 = ~n19583 & ~n19584;
  assign n19586 = ~n19582 & n19585;
  assign n19587 = n7294 & n12999;
  assign n19588 = n19586 & ~n19587;
  assign n19589 =  a[11]  & ~n19588;
  assign n19590 = ~n19588 & ~n19589;
  assign n19591 =  a[11]  & ~n19589;
  assign n19592 = ~n19590 & ~n19591;
  assign n19593 = ~n19448 & ~n19452;
  assign n19594 = ~n19451 & ~n19452;
  assign n19595 = ~n19593 & ~n19594;
  assign n19596 = ~n19592 & ~n19595;
  assign n19597 = ~n19592 & ~n19596;
  assign n19598 = ~n19595 & ~n19596;
  assign n19599 = ~n19597 & ~n19598;
  assign n19600 = n7983 & n12502;
  assign n19601 = n7291 & n12505;
  assign n19602 = n7632 & n12370;
  assign n19603 = ~n19601 & ~n19602;
  assign n19604 = ~n19600 & n19603;
  assign n19605 = n7294 & ~n13736;
  assign n19606 = n19604 & ~n19605;
  assign n19607 =  a[11]  & ~n19606;
  assign n19608 = ~n19606 & ~n19607;
  assign n19609 =  a[11]  & ~n19607;
  assign n19610 = ~n19608 & ~n19609;
  assign n19611 = ~n19443 & ~n19447;
  assign n19612 = ~n19446 & ~n19447;
  assign n19613 = ~n19611 & ~n19612;
  assign n19614 = ~n19610 & ~n19613;
  assign n19615 = ~n19610 & ~n19614;
  assign n19616 = ~n19613 & ~n19614;
  assign n19617 = ~n19615 & ~n19616;
  assign n19618 = n7983 & n12370;
  assign n19619 = n7291 & n12508;
  assign n19620 = n7632 & n12505;
  assign n19621 = ~n19619 & ~n19620;
  assign n19622 = ~n19618 & n19621;
  assign n19623 = n7294 & ~n13748;
  assign n19624 = n19622 & ~n19623;
  assign n19625 =  a[11]  & ~n19624;
  assign n19626 = ~n19624 & ~n19625;
  assign n19627 =  a[11]  & ~n19625;
  assign n19628 = ~n19626 & ~n19627;
  assign n19629 = ~n19438 & ~n19442;
  assign n19630 = ~n19441 & ~n19442;
  assign n19631 = ~n19629 & ~n19630;
  assign n19632 = ~n19628 & ~n19631;
  assign n19633 = ~n19628 & ~n19632;
  assign n19634 = ~n19631 & ~n19632;
  assign n19635 = ~n19633 & ~n19634;
  assign n19636 = n7983 & n12505;
  assign n19637 = n7291 & n12513;
  assign n19638 = n7632 & n12508;
  assign n19639 = ~n19637 & ~n19638;
  assign n19640 = ~n19636 & n19639;
  assign n19641 = n7294 & ~n14051;
  assign n19642 = n19640 & ~n19641;
  assign n19643 =  a[11]  & ~n19642;
  assign n19644 = ~n19642 & ~n19643;
  assign n19645 =  a[11]  & ~n19643;
  assign n19646 = ~n19644 & ~n19645;
  assign n19647 = ~n19433 & ~n19437;
  assign n19648 = ~n19436 & ~n19437;
  assign n19649 = ~n19647 & ~n19648;
  assign n19650 = ~n19646 & ~n19649;
  assign n19651 = ~n19646 & ~n19650;
  assign n19652 = ~n19649 & ~n19650;
  assign n19653 = ~n19651 & ~n19652;
  assign n19654 = n7983 & n12508;
  assign n19655 = n7291 & n12511;
  assign n19656 = n7632 & n12513;
  assign n19657 = ~n19655 & ~n19656;
  assign n19658 = ~n19654 & n19657;
  assign n19659 = n7294 & n13863;
  assign n19660 = n19658 & ~n19659;
  assign n19661 =  a[11]  & ~n19660;
  assign n19662 = ~n19660 & ~n19661;
  assign n19663 =  a[11]  & ~n19661;
  assign n19664 = ~n19662 & ~n19663;
  assign n19665 = ~n19428 & ~n19432;
  assign n19666 = ~n19431 & ~n19432;
  assign n19667 = ~n19665 & ~n19666;
  assign n19668 = ~n19664 & ~n19667;
  assign n19669 = ~n19664 & ~n19668;
  assign n19670 = ~n19667 & ~n19668;
  assign n19671 = ~n19669 & ~n19670;
  assign n19672 = n7983 & n12513;
  assign n19673 = n7291 & n12516;
  assign n19674 = n7632 & n12511;
  assign n19675 = ~n19673 & ~n19674;
  assign n19676 = ~n19672 & n19675;
  assign n19677 = n7294 & n14177;
  assign n19678 = n19676 & ~n19677;
  assign n19679 =  a[11]  & ~n19678;
  assign n19680 = ~n19678 & ~n19679;
  assign n19681 =  a[11]  & ~n19679;
  assign n19682 = ~n19680 & ~n19681;
  assign n19683 = ~n19423 & ~n19427;
  assign n19684 = ~n19426 & ~n19427;
  assign n19685 = ~n19683 & ~n19684;
  assign n19686 = ~n19682 & ~n19685;
  assign n19687 = ~n19682 & ~n19686;
  assign n19688 = ~n19685 & ~n19686;
  assign n19689 = ~n19687 & ~n19688;
  assign n19690 = n7983 & n12511;
  assign n19691 = n7291 & n12519;
  assign n19692 = n7632 & n12516;
  assign n19693 = ~n19691 & ~n19692;
  assign n19694 = ~n19690 & n19693;
  assign n19695 = n7294 & ~n14233;
  assign n19696 = n19694 & ~n19695;
  assign n19697 =  a[11]  & ~n19696;
  assign n19698 = ~n19696 & ~n19697;
  assign n19699 =  a[11]  & ~n19697;
  assign n19700 = ~n19698 & ~n19699;
  assign n19701 = ~n19418 & ~n19422;
  assign n19702 = ~n19421 & ~n19422;
  assign n19703 = ~n19701 & ~n19702;
  assign n19704 = ~n19700 & ~n19703;
  assign n19705 = ~n19700 & ~n19704;
  assign n19706 = ~n19703 & ~n19704;
  assign n19707 = ~n19705 & ~n19706;
  assign n19708 = n19109 & n19416;
  assign n19709 = ~n19417 & ~n19708;
  assign n19710 = n7983 & n12516;
  assign n19711 = n7291 & n12522;
  assign n19712 = n7632 & n12519;
  assign n19713 = ~n19711 & ~n19712;
  assign n19714 = ~n19710 & n19713;
  assign n19715 = ~n7294 & n19714;
  assign n19716 = n14443 & n19714;
  assign n19717 = ~n19715 & ~n19716;
  assign n19718 =  a[11]  & ~n19717;
  assign n19719 = ~ a[11]  & n19717;
  assign n19720 = ~n19718 & ~n19719;
  assign n19721 = n19709 & ~n19720;
  assign n19722 = n19127 & n19414;
  assign n19723 = ~n19415 & ~n19722;
  assign n19724 = n7983 & n12519;
  assign n19725 = n7291 & n12525;
  assign n19726 = n7632 & n12522;
  assign n19727 = ~n19725 & ~n19726;
  assign n19728 = ~n19724 & n19727;
  assign n19729 = ~n7294 & n19728;
  assign n19730 = ~n14454 & n19728;
  assign n19731 = ~n19729 & ~n19730;
  assign n19732 =  a[11]  & ~n19731;
  assign n19733 = ~ a[11]  & n19731;
  assign n19734 = ~n19732 & ~n19733;
  assign n19735 = n19723 & ~n19734;
  assign n19736 = n7983 & n12522;
  assign n19737 = n7291 & n12528;
  assign n19738 = n7632 & n12525;
  assign n19739 = ~n19737 & ~n19738;
  assign n19740 = ~n19736 & n19739;
  assign n19741 = n7294 & n14837;
  assign n19742 = n19740 & ~n19741;
  assign n19743 =  a[11]  & ~n19742;
  assign n19744 = ~n19742 & ~n19743;
  assign n19745 =  a[11]  & ~n19743;
  assign n19746 = ~n19744 & ~n19745;
  assign n19747 = n19410 & ~n19412;
  assign n19748 = ~n19413 & ~n19747;
  assign n19749 = ~n19746 & n19748;
  assign n19750 = ~n19746 & ~n19749;
  assign n19751 = n19748 & ~n19749;
  assign n19752 = ~n19750 & ~n19751;
  assign n19753 = n7983 & n12525;
  assign n19754 = n7291 & n12531;
  assign n19755 = n7632 & n12528;
  assign n19756 = ~n19754 & ~n19755;
  assign n19757 = ~n19753 & n19756;
  assign n19758 = n7294 & n14608;
  assign n19759 = n19757 & ~n19758;
  assign n19760 =  a[11]  & ~n19759;
  assign n19761 = ~n19759 & ~n19760;
  assign n19762 =  a[11]  & ~n19760;
  assign n19763 = ~n19761 & ~n19762;
  assign n19764 = ~n19405 & ~n19409;
  assign n19765 = ~n19408 & ~n19409;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~n19763 & ~n19766;
  assign n19768 = ~n19763 & ~n19767;
  assign n19769 = ~n19766 & ~n19767;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = n7983 & n12528;
  assign n19772 = n7291 & n12534;
  assign n19773 = n7632 & n12531;
  assign n19774 = ~n19772 & ~n19773;
  assign n19775 = ~n19771 & n19774;
  assign n19776 = n7294 & ~n15003;
  assign n19777 = n19775 & ~n19776;
  assign n19778 =  a[11]  & ~n19777;
  assign n19779 = ~n19777 & ~n19778;
  assign n19780 =  a[11]  & ~n19778;
  assign n19781 = ~n19779 & ~n19780;
  assign n19782 = ~n19400 & ~n19404;
  assign n19783 = ~n19403 & ~n19404;
  assign n19784 = ~n19782 & ~n19783;
  assign n19785 = ~n19781 & ~n19784;
  assign n19786 = ~n19781 & ~n19785;
  assign n19787 = ~n19784 & ~n19785;
  assign n19788 = ~n19786 & ~n19787;
  assign n19789 = n19186 & n19398;
  assign n19790 = ~n19399 & ~n19789;
  assign n19791 = n7983 & n12531;
  assign n19792 = n7291 & n12537;
  assign n19793 = n7632 & n12534;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = ~n19791 & n19794;
  assign n19796 = ~n7294 & n19795;
  assign n19797 = ~n15255 & n19795;
  assign n19798 = ~n19796 & ~n19797;
  assign n19799 =  a[11]  & ~n19798;
  assign n19800 = ~ a[11]  & n19798;
  assign n19801 = ~n19799 & ~n19800;
  assign n19802 = n19790 & ~n19801;
  assign n19803 = n19204 & n19396;
  assign n19804 = ~n19397 & ~n19803;
  assign n19805 = n7983 & n12534;
  assign n19806 = n7291 & n12540;
  assign n19807 = n7632 & n12537;
  assign n19808 = ~n19806 & ~n19807;
  assign n19809 = ~n19805 & n19808;
  assign n19810 = ~n7294 & n19809;
  assign n19811 = n15096 & n19809;
  assign n19812 = ~n19810 & ~n19811;
  assign n19813 =  a[11]  & ~n19812;
  assign n19814 = ~ a[11]  & n19812;
  assign n19815 = ~n19813 & ~n19814;
  assign n19816 = n19804 & ~n19815;
  assign n19817 = n19222 & n19394;
  assign n19818 = ~n19395 & ~n19817;
  assign n19819 = n7983 & n12537;
  assign n19820 = n7291 & n12543;
  assign n19821 = n7632 & n12540;
  assign n19822 = ~n19820 & ~n19821;
  assign n19823 = ~n19819 & n19822;
  assign n19824 = ~n7294 & n19823;
  assign n19825 = n15385 & n19823;
  assign n19826 = ~n19824 & ~n19825;
  assign n19827 =  a[11]  & ~n19826;
  assign n19828 = ~ a[11]  & n19826;
  assign n19829 = ~n19827 & ~n19828;
  assign n19830 = n19818 & ~n19829;
  assign n19831 = n7983 & n12540;
  assign n19832 = n7291 & n12546;
  assign n19833 = n7632 & n12543;
  assign n19834 = ~n19832 & ~n19833;
  assign n19835 = ~n19831 & n19834;
  assign n19836 = n7294 & ~n15708;
  assign n19837 = n19835 & ~n19836;
  assign n19838 =  a[11]  & ~n19837;
  assign n19839 = ~n19837 & ~n19838;
  assign n19840 =  a[11]  & ~n19838;
  assign n19841 = ~n19839 & ~n19840;
  assign n19842 = n19390 & ~n19392;
  assign n19843 = ~n19393 & ~n19842;
  assign n19844 = ~n19841 & n19843;
  assign n19845 = ~n19841 & ~n19844;
  assign n19846 = n19843 & ~n19844;
  assign n19847 = ~n19845 & ~n19846;
  assign n19848 = n7983 & n12543;
  assign n19849 = n7291 & n12549;
  assign n19850 = n7632 & n12546;
  assign n19851 = ~n19849 & ~n19850;
  assign n19852 = ~n19848 & n19851;
  assign n19853 = n7294 & n15724;
  assign n19854 = n19852 & ~n19853;
  assign n19855 =  a[11]  & ~n19854;
  assign n19856 = ~n19854 & ~n19855;
  assign n19857 =  a[11]  & ~n19855;
  assign n19858 = ~n19856 & ~n19857;
  assign n19859 = ~n19385 & ~n19389;
  assign n19860 = ~n19388 & ~n19389;
  assign n19861 = ~n19859 & ~n19860;
  assign n19862 = ~n19858 & ~n19861;
  assign n19863 = ~n19858 & ~n19862;
  assign n19864 = ~n19861 & ~n19862;
  assign n19865 = ~n19863 & ~n19864;
  assign n19866 = n7983 & n12546;
  assign n19867 = n7291 & n12552;
  assign n19868 = n7632 & n12549;
  assign n19869 = ~n19867 & ~n19868;
  assign n19870 = ~n19866 & n19869;
  assign n19871 = n7294 & ~n15356;
  assign n19872 = n19870 & ~n19871;
  assign n19873 =  a[11]  & ~n19872;
  assign n19874 = ~n19872 & ~n19873;
  assign n19875 =  a[11]  & ~n19873;
  assign n19876 = ~n19874 & ~n19875;
  assign n19877 = ~n19380 & ~n19384;
  assign n19878 = ~n19383 & ~n19384;
  assign n19879 = ~n19877 & ~n19878;
  assign n19880 = ~n19876 & ~n19879;
  assign n19881 = ~n19876 & ~n19880;
  assign n19882 = ~n19879 & ~n19880;
  assign n19883 = ~n19881 & ~n19882;
  assign n19884 = n19281 & n19378;
  assign n19885 = ~n19379 & ~n19884;
  assign n19886 = n7983 & n12549;
  assign n19887 = n7291 & n12555;
  assign n19888 = n7632 & n12552;
  assign n19889 = ~n19887 & ~n19888;
  assign n19890 = ~n19886 & n19889;
  assign n19891 = ~n7294 & n19890;
  assign n19892 = ~n15764 & n19890;
  assign n19893 = ~n19891 & ~n19892;
  assign n19894 =  a[11]  & ~n19893;
  assign n19895 = ~ a[11]  & n19893;
  assign n19896 = ~n19894 & ~n19895;
  assign n19897 = n19885 & ~n19896;
  assign n19898 = n19374 & ~n19376;
  assign n19899 = ~n19377 & ~n19898;
  assign n19900 = n7983 & n12552;
  assign n19901 = n7291 & n12558;
  assign n19902 = n7632 & n12555;
  assign n19903 = ~n19901 & ~n19902;
  assign n19904 = ~n19900 & n19903;
  assign n19905 = ~n7294 & n19904;
  assign n19906 = n15791 & n19904;
  assign n19907 = ~n19905 & ~n19906;
  assign n19908 =  a[11]  & ~n19907;
  assign n19909 = ~ a[11]  & n19907;
  assign n19910 = ~n19908 & ~n19909;
  assign n19911 = n19899 & ~n19910;
  assign n19912 = n19313 & n19372;
  assign n19913 = ~n19373 & ~n19912;
  assign n19914 = n7983 & n12555;
  assign n19915 = n7291 & n12561;
  assign n19916 = n7632 & n12558;
  assign n19917 = ~n19915 & ~n19916;
  assign n19918 = ~n19914 & n19917;
  assign n19919 = ~n7294 & n19918;
  assign n19920 = n15816 & n19918;
  assign n19921 = ~n19919 & ~n19920;
  assign n19922 =  a[11]  & ~n19921;
  assign n19923 = ~ a[11]  & n19921;
  assign n19924 = ~n19922 & ~n19923;
  assign n19925 = n19913 & ~n19924;
  assign n19926 = n7983 & n12558;
  assign n19927 = n7291 & n12564;
  assign n19928 = n7632 & n12561;
  assign n19929 = ~n19927 & ~n19928;
  assign n19930 = ~n19926 & n19929;
  assign n19931 = n7294 & n15847;
  assign n19932 = n19930 & ~n19931;
  assign n19933 =  a[11]  & ~n19932;
  assign n19934 = ~n19932 & ~n19933;
  assign n19935 =  a[11]  & ~n19933;
  assign n19936 = ~n19934 & ~n19935;
  assign n19937 = n19368 & ~n19370;
  assign n19938 = ~n19371 & ~n19937;
  assign n19939 = ~n19936 & n19938;
  assign n19940 = ~n19936 & ~n19939;
  assign n19941 = n19938 & ~n19939;
  assign n19942 = ~n19940 & ~n19941;
  assign n19943 = ~n19355 & ~n19367;
  assign n19944 = ~n19366 & ~n19367;
  assign n19945 = ~n19943 & ~n19944;
  assign n19946 = n7983 & n12561;
  assign n19947 = n7291 & n12567;
  assign n19948 = n7632 & n12564;
  assign n19949 = ~n19947 & ~n19948;
  assign n19950 = ~n19946 & n19949;
  assign n19951 = ~n7294 & n19950;
  assign n19952 = n15905 & n19950;
  assign n19953 = ~n19951 & ~n19952;
  assign n19954 =  a[11]  & ~n19953;
  assign n19955 = ~ a[11]  & n19953;
  assign n19956 = ~n19954 & ~n19955;
  assign n19957 = ~n19945 & ~n19956;
  assign n19958 = n7983 & n12564;
  assign n19959 = n7291 & n12571;
  assign n19960 = n7632 & n12567;
  assign n19961 = ~n19959 & ~n19960;
  assign n19962 = ~n19958 & n19961;
  assign n19963 = n7294 & ~n15944;
  assign n19964 = n19962 & ~n19963;
  assign n19965 =  a[11]  & ~n19964;
  assign n19966 = ~n19964 & ~n19965;
  assign n19967 =  a[11]  & ~n19965;
  assign n19968 = ~n19966 & ~n19967;
  assign n19969 = ~n19339 & n19350;
  assign n19970 = ~n19351 & ~n19969;
  assign n19971 = ~n19968 & n19970;
  assign n19972 = ~n19968 & ~n19971;
  assign n19973 = n19970 & ~n19971;
  assign n19974 = ~n19972 & ~n19973;
  assign n19975 = n19336 & ~n19338;
  assign n19976 = ~n19339 & ~n19975;
  assign n19977 = n7983 & n12567;
  assign n19978 = n7291 & n12574;
  assign n19979 = n7632 & n12571;
  assign n19980 = ~n19978 & ~n19979;
  assign n19981 = ~n19977 & n19980;
  assign n19982 = ~n7294 & n19981;
  assign n19983 = ~n15989 & n19981;
  assign n19984 = ~n19982 & ~n19983;
  assign n19985 =  a[11]  & ~n19984;
  assign n19986 = ~ a[11]  & n19984;
  assign n19987 = ~n19985 & ~n19986;
  assign n19988 = n19976 & ~n19987;
  assign n19989 = n7632 & ~n12581;
  assign n19990 = n7983 & n12577;
  assign n19991 = ~n19989 & ~n19990;
  assign n19992 = n7294 & ~n16085;
  assign n19993 = n19991 & ~n19992;
  assign n19994 =  a[11]  & ~n19993;
  assign n19995 =  a[11]  & ~n19994;
  assign n19996 = ~n19993 & ~n19994;
  assign n19997 = ~n19995 & ~n19996;
  assign n19998 = ~n7289 & ~n12581;
  assign n19999 =  a[11]  & ~n19998;
  assign n20000 = ~n19997 & n19999;
  assign n20001 = n7983 & n12574;
  assign n20002 = n7291 & ~n12581;
  assign n20003 = n7632 & n12577;
  assign n20004 = ~n20002 & ~n20003;
  assign n20005 = ~n20001 & n20004;
  assign n20006 = ~n7294 & n20005;
  assign n20007 = n16094 & n20005;
  assign n20008 = ~n20006 & ~n20007;
  assign n20009 =  a[11]  & ~n20008;
  assign n20010 = ~ a[11]  & n20008;
  assign n20011 = ~n20009 & ~n20010;
  assign n20012 = n20000 & ~n20011;
  assign n20013 = n19337 & n20012;
  assign n20014 = n20012 & ~n20013;
  assign n20015 = n19337 & ~n20013;
  assign n20016 = ~n20014 & ~n20015;
  assign n20017 = n7983 & n12571;
  assign n20018 = n7291 & n12577;
  assign n20019 = n7632 & n12574;
  assign n20020 = ~n20018 & ~n20019;
  assign n20021 = ~n20017 & n20020;
  assign n20022 = n7294 & n16013;
  assign n20023 = n20021 & ~n20022;
  assign n20024 =  a[11]  & ~n20023;
  assign n20025 =  a[11]  & ~n20024;
  assign n20026 = ~n20023 & ~n20024;
  assign n20027 = ~n20025 & ~n20026;
  assign n20028 = ~n20016 & ~n20027;
  assign n20029 = ~n20013 & ~n20028;
  assign n20030 = ~n19976 & n19987;
  assign n20031 = ~n19988 & ~n20030;
  assign n20032 = ~n20029 & n20031;
  assign n20033 = ~n19988 & ~n20032;
  assign n20034 = ~n19974 & ~n20033;
  assign n20035 = ~n19971 & ~n20034;
  assign n20036 = n19945 & n19956;
  assign n20037 = ~n19957 & ~n20036;
  assign n20038 = ~n20035 & n20037;
  assign n20039 = ~n19957 & ~n20038;
  assign n20040 = ~n19942 & ~n20039;
  assign n20041 = ~n19939 & ~n20040;
  assign n20042 = n19913 & ~n19925;
  assign n20043 = ~n19924 & ~n19925;
  assign n20044 = ~n20042 & ~n20043;
  assign n20045 = ~n20041 & ~n20044;
  assign n20046 = ~n19925 & ~n20045;
  assign n20047 = n19899 & ~n19911;
  assign n20048 = ~n19910 & ~n19911;
  assign n20049 = ~n20047 & ~n20048;
  assign n20050 = ~n20046 & ~n20049;
  assign n20051 = ~n19911 & ~n20050;
  assign n20052 = ~n19885 & n19896;
  assign n20053 = ~n19897 & ~n20052;
  assign n20054 = ~n20051 & n20053;
  assign n20055 = ~n19897 & ~n20054;
  assign n20056 = ~n19883 & ~n20055;
  assign n20057 = ~n19880 & ~n20056;
  assign n20058 = ~n19865 & ~n20057;
  assign n20059 = ~n19862 & ~n20058;
  assign n20060 = ~n19847 & ~n20059;
  assign n20061 = ~n19844 & ~n20060;
  assign n20062 = n19818 & ~n19830;
  assign n20063 = ~n19829 & ~n19830;
  assign n20064 = ~n20062 & ~n20063;
  assign n20065 = ~n20061 & ~n20064;
  assign n20066 = ~n19830 & ~n20065;
  assign n20067 = n19804 & ~n19816;
  assign n20068 = ~n19815 & ~n19816;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = ~n20066 & ~n20069;
  assign n20071 = ~n19816 & ~n20070;
  assign n20072 = ~n19790 & n19801;
  assign n20073 = ~n19802 & ~n20072;
  assign n20074 = ~n20071 & n20073;
  assign n20075 = ~n19802 & ~n20074;
  assign n20076 = ~n19788 & ~n20075;
  assign n20077 = ~n19785 & ~n20076;
  assign n20078 = ~n19770 & ~n20077;
  assign n20079 = ~n19767 & ~n20078;
  assign n20080 = ~n19752 & ~n20079;
  assign n20081 = ~n19749 & ~n20080;
  assign n20082 = n19723 & ~n19735;
  assign n20083 = ~n19734 & ~n19735;
  assign n20084 = ~n20082 & ~n20083;
  assign n20085 = ~n20081 & ~n20084;
  assign n20086 = ~n19735 & ~n20085;
  assign n20087 = ~n19709 & n19720;
  assign n20088 = ~n19721 & ~n20087;
  assign n20089 = ~n20086 & n20088;
  assign n20090 = ~n19721 & ~n20089;
  assign n20091 = ~n19707 & ~n20090;
  assign n20092 = ~n19704 & ~n20091;
  assign n20093 = ~n19689 & ~n20092;
  assign n20094 = ~n19686 & ~n20093;
  assign n20095 = ~n19671 & ~n20094;
  assign n20096 = ~n19668 & ~n20095;
  assign n20097 = ~n19653 & ~n20096;
  assign n20098 = ~n19650 & ~n20097;
  assign n20099 = ~n19635 & ~n20098;
  assign n20100 = ~n19632 & ~n20099;
  assign n20101 = ~n19617 & ~n20100;
  assign n20102 = ~n19614 & ~n20101;
  assign n20103 = ~n19599 & ~n20102;
  assign n20104 = ~n19596 & ~n20103;
  assign n20105 = ~n19581 & ~n20104;
  assign n20106 = ~n19578 & ~n20105;
  assign n20107 = ~n19563 & ~n20106;
  assign n20108 = ~n19560 & ~n20107;
  assign n20109 = ~n19545 & ~n20108;
  assign n20110 = ~n19542 & ~n20109;
  assign n20111 = ~n19528 & ~n20110;
  assign n20112 = n19528 & n20110;
  assign n20113 = ~n20111 & ~n20112;
  assign n20114 = n9331 & n13630;
  assign n20115 = n8418 & n13515;
  assign n20116 = n8860 & n13597;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = ~n20114 & n20117;
  assign n20119 = n8421 & n13976;
  assign n20120 = n20118 & ~n20119;
  assign n20121 =  a[8]  & ~n20120;
  assign n20122 =  a[8]  & ~n20121;
  assign n20123 = ~n20120 & ~n20121;
  assign n20124 = ~n20122 & ~n20123;
  assign n20125 = n20113 & ~n20124;
  assign n20126 = ~n20111 & ~n20125;
  assign n20127 = ~n19525 & ~n20126;
  assign n20128 = n19525 & n20126;
  assign n20129 = ~n20127 & ~n20128;
  assign n20130 = n71 & ~n13438;
  assign n20131 = n9867 & ~n13627;
  assign n20132 = n10434 & n13941;
  assign n20133 = ~n20131 & ~n20132;
  assign n20134 = ~n20130 & n20133;
  assign n20135 = n9870 & n14028;
  assign n20136 = n20134 & ~n20135;
  assign n20137 =  a[5]  & ~n20136;
  assign n20138 =  a[5]  & ~n20137;
  assign n20139 = ~n20136 & ~n20137;
  assign n20140 = ~n20138 & ~n20139;
  assign n20141 = n20129 & ~n20140;
  assign n20142 = ~n20127 & ~n20141;
  assign n20143 = ~n19522 & ~n20142;
  assign n20144 = n19522 & n20142;
  assign n20145 = ~n20143 & ~n20144;
  assign n20146 = n20129 & ~n20141;
  assign n20147 = ~n20140 & ~n20141;
  assign n20148 = ~n20146 & ~n20147;
  assign n20149 = n20113 & ~n20125;
  assign n20150 = ~n20124 & ~n20125;
  assign n20151 = ~n20149 & ~n20150;
  assign n20152 = n19545 & n20108;
  assign n20153 = ~n20109 & ~n20152;
  assign n20154 = n9331 & n13597;
  assign n20155 = n8418 & n13521;
  assign n20156 = n8860 & n13515;
  assign n20157 = ~n20155 & ~n20156;
  assign n20158 = ~n20154 & n20157;
  assign n20159 = ~n8421 & n20158;
  assign n20160 = n13612 & n20158;
  assign n20161 = ~n20159 & ~n20160;
  assign n20162 =  a[8]  & ~n20161;
  assign n20163 = ~ a[8]  & n20161;
  assign n20164 = ~n20162 & ~n20163;
  assign n20165 = n20153 & ~n20164;
  assign n20166 = n19563 & n20106;
  assign n20167 = ~n20107 & ~n20166;
  assign n20168 = n9331 & n13515;
  assign n20169 = n8418 & n13518;
  assign n20170 = n8860 & n13521;
  assign n20171 = ~n20169 & ~n20170;
  assign n20172 = ~n20168 & n20171;
  assign n20173 = ~n8421 & n20172;
  assign n20174 = ~n13541 & n20172;
  assign n20175 = ~n20173 & ~n20174;
  assign n20176 =  a[8]  & ~n20175;
  assign n20177 = ~ a[8]  & n20175;
  assign n20178 = ~n20176 & ~n20177;
  assign n20179 = n20167 & ~n20178;
  assign n20180 = n19581 & n20104;
  assign n20181 = ~n20105 & ~n20180;
  assign n20182 = n9331 & n13521;
  assign n20183 = n8418 & n13491;
  assign n20184 = n8860 & n13518;
  assign n20185 = ~n20183 & ~n20184;
  assign n20186 = ~n20182 & n20185;
  assign n20187 = ~n8421 & n20186;
  assign n20188 = n13909 & n20186;
  assign n20189 = ~n20187 & ~n20188;
  assign n20190 =  a[8]  & ~n20189;
  assign n20191 = ~ a[8]  & n20189;
  assign n20192 = ~n20190 & ~n20191;
  assign n20193 = n20181 & ~n20192;
  assign n20194 = n19599 & n20102;
  assign n20195 = ~n20103 & ~n20194;
  assign n20196 = n9331 & n13518;
  assign n20197 = n8418 & n12889;
  assign n20198 = n8860 & n13491;
  assign n20199 = ~n20197 & ~n20198;
  assign n20200 = ~n20196 & n20199;
  assign n20201 = ~n8421 & n20200;
  assign n20202 = ~n13584 & n20200;
  assign n20203 = ~n20201 & ~n20202;
  assign n20204 =  a[8]  & ~n20203;
  assign n20205 = ~ a[8]  & n20203;
  assign n20206 = ~n20204 & ~n20205;
  assign n20207 = n20195 & ~n20206;
  assign n20208 = n19617 & n20100;
  assign n20209 = ~n20101 & ~n20208;
  assign n20210 = n9331 & n13491;
  assign n20211 = n8418 & n12769;
  assign n20212 = n8860 & n12889;
  assign n20213 = ~n20211 & ~n20212;
  assign n20214 = ~n20210 & n20213;
  assign n20215 = ~n8421 & n20214;
  assign n20216 = n13503 & n20214;
  assign n20217 = ~n20215 & ~n20216;
  assign n20218 =  a[8]  & ~n20217;
  assign n20219 = ~ a[8]  & n20217;
  assign n20220 = ~n20218 & ~n20219;
  assign n20221 = n20209 & ~n20220;
  assign n20222 = n19635 & n20098;
  assign n20223 = ~n20099 & ~n20222;
  assign n20224 = n9331 & n12889;
  assign n20225 = n8418 & n12502;
  assign n20226 = n8860 & n12769;
  assign n20227 = ~n20225 & ~n20226;
  assign n20228 = ~n20224 & n20227;
  assign n20229 = ~n8421 & n20228;
  assign n20230 = ~n12895 & n20228;
  assign n20231 = ~n20229 & ~n20230;
  assign n20232 =  a[8]  & ~n20231;
  assign n20233 = ~ a[8]  & n20231;
  assign n20234 = ~n20232 & ~n20233;
  assign n20235 = n20223 & ~n20234;
  assign n20236 = n19653 & n20096;
  assign n20237 = ~n20097 & ~n20236;
  assign n20238 = n9331 & n12769;
  assign n20239 = n8418 & n12370;
  assign n20240 = n8860 & n12502;
  assign n20241 = ~n20239 & ~n20240;
  assign n20242 = ~n20238 & n20241;
  assign n20243 = ~n8421 & n20242;
  assign n20244 = ~n12999 & n20242;
  assign n20245 = ~n20243 & ~n20244;
  assign n20246 =  a[8]  & ~n20245;
  assign n20247 = ~ a[8]  & n20245;
  assign n20248 = ~n20246 & ~n20247;
  assign n20249 = n20237 & ~n20248;
  assign n20250 = n19671 & n20094;
  assign n20251 = ~n20095 & ~n20250;
  assign n20252 = n9331 & n12502;
  assign n20253 = n8418 & n12505;
  assign n20254 = n8860 & n12370;
  assign n20255 = ~n20253 & ~n20254;
  assign n20256 = ~n20252 & n20255;
  assign n20257 = ~n8421 & n20256;
  assign n20258 = n13736 & n20256;
  assign n20259 = ~n20257 & ~n20258;
  assign n20260 =  a[8]  & ~n20259;
  assign n20261 = ~ a[8]  & n20259;
  assign n20262 = ~n20260 & ~n20261;
  assign n20263 = n20251 & ~n20262;
  assign n20264 = n19689 & n20092;
  assign n20265 = ~n20093 & ~n20264;
  assign n20266 = n9331 & n12370;
  assign n20267 = n8418 & n12508;
  assign n20268 = n8860 & n12505;
  assign n20269 = ~n20267 & ~n20268;
  assign n20270 = ~n20266 & n20269;
  assign n20271 = ~n8421 & n20270;
  assign n20272 = n13748 & n20270;
  assign n20273 = ~n20271 & ~n20272;
  assign n20274 =  a[8]  & ~n20273;
  assign n20275 = ~ a[8]  & n20273;
  assign n20276 = ~n20274 & ~n20275;
  assign n20277 = n20265 & ~n20276;
  assign n20278 = n19707 & n20090;
  assign n20279 = ~n20091 & ~n20278;
  assign n20280 = n9331 & n12505;
  assign n20281 = n8418 & n12513;
  assign n20282 = n8860 & n12508;
  assign n20283 = ~n20281 & ~n20282;
  assign n20284 = ~n20280 & n20283;
  assign n20285 = ~n8421 & n20284;
  assign n20286 = n14051 & n20284;
  assign n20287 = ~n20285 & ~n20286;
  assign n20288 =  a[8]  & ~n20287;
  assign n20289 = ~ a[8]  & n20287;
  assign n20290 = ~n20288 & ~n20289;
  assign n20291 = n20279 & ~n20290;
  assign n20292 = n9331 & n12508;
  assign n20293 = n8418 & n12511;
  assign n20294 = n8860 & n12513;
  assign n20295 = ~n20293 & ~n20294;
  assign n20296 = ~n20292 & n20295;
  assign n20297 = n8421 & n13863;
  assign n20298 = n20296 & ~n20297;
  assign n20299 =  a[8]  & ~n20298;
  assign n20300 = ~n20298 & ~n20299;
  assign n20301 =  a[8]  & ~n20299;
  assign n20302 = ~n20300 & ~n20301;
  assign n20303 = n20086 & ~n20088;
  assign n20304 = ~n20089 & ~n20303;
  assign n20305 = ~n20302 & n20304;
  assign n20306 = ~n20302 & ~n20305;
  assign n20307 = n20304 & ~n20305;
  assign n20308 = ~n20306 & ~n20307;
  assign n20309 = n9331 & n12513;
  assign n20310 = n8418 & n12516;
  assign n20311 = n8860 & n12511;
  assign n20312 = ~n20310 & ~n20311;
  assign n20313 = ~n20309 & n20312;
  assign n20314 = n8421 & n14177;
  assign n20315 = n20313 & ~n20314;
  assign n20316 =  a[8]  & ~n20315;
  assign n20317 = ~n20315 & ~n20316;
  assign n20318 =  a[8]  & ~n20316;
  assign n20319 = ~n20317 & ~n20318;
  assign n20320 = ~n20081 & ~n20085;
  assign n20321 = ~n20084 & ~n20085;
  assign n20322 = ~n20320 & ~n20321;
  assign n20323 = ~n20319 & ~n20322;
  assign n20324 = ~n20319 & ~n20323;
  assign n20325 = ~n20322 & ~n20323;
  assign n20326 = ~n20324 & ~n20325;
  assign n20327 = n19752 & n20079;
  assign n20328 = ~n20080 & ~n20327;
  assign n20329 = n9331 & n12511;
  assign n20330 = n8418 & n12519;
  assign n20331 = n8860 & n12516;
  assign n20332 = ~n20330 & ~n20331;
  assign n20333 = ~n20329 & n20332;
  assign n20334 = ~n8421 & n20333;
  assign n20335 = n14233 & n20333;
  assign n20336 = ~n20334 & ~n20335;
  assign n20337 =  a[8]  & ~n20336;
  assign n20338 = ~ a[8]  & n20336;
  assign n20339 = ~n20337 & ~n20338;
  assign n20340 = n20328 & ~n20339;
  assign n20341 = n19770 & n20077;
  assign n20342 = ~n20078 & ~n20341;
  assign n20343 = n9331 & n12516;
  assign n20344 = n8418 & n12522;
  assign n20345 = n8860 & n12519;
  assign n20346 = ~n20344 & ~n20345;
  assign n20347 = ~n20343 & n20346;
  assign n20348 = ~n8421 & n20347;
  assign n20349 = n14443 & n20347;
  assign n20350 = ~n20348 & ~n20349;
  assign n20351 =  a[8]  & ~n20350;
  assign n20352 = ~ a[8]  & n20350;
  assign n20353 = ~n20351 & ~n20352;
  assign n20354 = n20342 & ~n20353;
  assign n20355 = n19788 & n20075;
  assign n20356 = ~n20076 & ~n20355;
  assign n20357 = n9331 & n12519;
  assign n20358 = n8418 & n12525;
  assign n20359 = n8860 & n12522;
  assign n20360 = ~n20358 & ~n20359;
  assign n20361 = ~n20357 & n20360;
  assign n20362 = ~n8421 & n20361;
  assign n20363 = ~n14454 & n20361;
  assign n20364 = ~n20362 & ~n20363;
  assign n20365 =  a[8]  & ~n20364;
  assign n20366 = ~ a[8]  & n20364;
  assign n20367 = ~n20365 & ~n20366;
  assign n20368 = n20356 & ~n20367;
  assign n20369 = n9331 & n12522;
  assign n20370 = n8418 & n12528;
  assign n20371 = n8860 & n12525;
  assign n20372 = ~n20370 & ~n20371;
  assign n20373 = ~n20369 & n20372;
  assign n20374 = n8421 & n14837;
  assign n20375 = n20373 & ~n20374;
  assign n20376 =  a[8]  & ~n20375;
  assign n20377 = ~n20375 & ~n20376;
  assign n20378 =  a[8]  & ~n20376;
  assign n20379 = ~n20377 & ~n20378;
  assign n20380 = n20071 & ~n20073;
  assign n20381 = ~n20074 & ~n20380;
  assign n20382 = ~n20379 & n20381;
  assign n20383 = ~n20379 & ~n20382;
  assign n20384 = n20381 & ~n20382;
  assign n20385 = ~n20383 & ~n20384;
  assign n20386 = n9331 & n12525;
  assign n20387 = n8418 & n12531;
  assign n20388 = n8860 & n12528;
  assign n20389 = ~n20387 & ~n20388;
  assign n20390 = ~n20386 & n20389;
  assign n20391 = n8421 & n14608;
  assign n20392 = n20390 & ~n20391;
  assign n20393 =  a[8]  & ~n20392;
  assign n20394 = ~n20392 & ~n20393;
  assign n20395 =  a[8]  & ~n20393;
  assign n20396 = ~n20394 & ~n20395;
  assign n20397 = ~n20066 & ~n20070;
  assign n20398 = ~n20069 & ~n20070;
  assign n20399 = ~n20397 & ~n20398;
  assign n20400 = ~n20396 & ~n20399;
  assign n20401 = ~n20396 & ~n20400;
  assign n20402 = ~n20399 & ~n20400;
  assign n20403 = ~n20401 & ~n20402;
  assign n20404 = n9331 & n12528;
  assign n20405 = n8418 & n12534;
  assign n20406 = n8860 & n12531;
  assign n20407 = ~n20405 & ~n20406;
  assign n20408 = ~n20404 & n20407;
  assign n20409 = n8421 & ~n15003;
  assign n20410 = n20408 & ~n20409;
  assign n20411 =  a[8]  & ~n20410;
  assign n20412 = ~n20410 & ~n20411;
  assign n20413 =  a[8]  & ~n20411;
  assign n20414 = ~n20412 & ~n20413;
  assign n20415 = ~n20061 & ~n20065;
  assign n20416 = ~n20064 & ~n20065;
  assign n20417 = ~n20415 & ~n20416;
  assign n20418 = ~n20414 & ~n20417;
  assign n20419 = ~n20414 & ~n20418;
  assign n20420 = ~n20417 & ~n20418;
  assign n20421 = ~n20419 & ~n20420;
  assign n20422 = n19847 & n20059;
  assign n20423 = ~n20060 & ~n20422;
  assign n20424 = n9331 & n12531;
  assign n20425 = n8418 & n12537;
  assign n20426 = n8860 & n12534;
  assign n20427 = ~n20425 & ~n20426;
  assign n20428 = ~n20424 & n20427;
  assign n20429 = ~n8421 & n20428;
  assign n20430 = ~n15255 & n20428;
  assign n20431 = ~n20429 & ~n20430;
  assign n20432 =  a[8]  & ~n20431;
  assign n20433 = ~ a[8]  & n20431;
  assign n20434 = ~n20432 & ~n20433;
  assign n20435 = n20423 & ~n20434;
  assign n20436 = n19865 & n20057;
  assign n20437 = ~n20058 & ~n20436;
  assign n20438 = n9331 & n12534;
  assign n20439 = n8418 & n12540;
  assign n20440 = n8860 & n12537;
  assign n20441 = ~n20439 & ~n20440;
  assign n20442 = ~n20438 & n20441;
  assign n20443 = ~n8421 & n20442;
  assign n20444 = n15096 & n20442;
  assign n20445 = ~n20443 & ~n20444;
  assign n20446 =  a[8]  & ~n20445;
  assign n20447 = ~ a[8]  & n20445;
  assign n20448 = ~n20446 & ~n20447;
  assign n20449 = n20437 & ~n20448;
  assign n20450 = n19883 & n20055;
  assign n20451 = ~n20056 & ~n20450;
  assign n20452 = n9331 & n12537;
  assign n20453 = n8418 & n12543;
  assign n20454 = n8860 & n12540;
  assign n20455 = ~n20453 & ~n20454;
  assign n20456 = ~n20452 & n20455;
  assign n20457 = ~n8421 & n20456;
  assign n20458 = n15385 & n20456;
  assign n20459 = ~n20457 & ~n20458;
  assign n20460 =  a[8]  & ~n20459;
  assign n20461 = ~ a[8]  & n20459;
  assign n20462 = ~n20460 & ~n20461;
  assign n20463 = n20451 & ~n20462;
  assign n20464 = n9331 & n12540;
  assign n20465 = n8418 & n12546;
  assign n20466 = n8860 & n12543;
  assign n20467 = ~n20465 & ~n20466;
  assign n20468 = ~n20464 & n20467;
  assign n20469 = n8421 & ~n15708;
  assign n20470 = n20468 & ~n20469;
  assign n20471 =  a[8]  & ~n20470;
  assign n20472 = ~n20470 & ~n20471;
  assign n20473 =  a[8]  & ~n20471;
  assign n20474 = ~n20472 & ~n20473;
  assign n20475 = n20051 & ~n20053;
  assign n20476 = ~n20054 & ~n20475;
  assign n20477 = ~n20474 & n20476;
  assign n20478 = ~n20474 & ~n20477;
  assign n20479 = n20476 & ~n20477;
  assign n20480 = ~n20478 & ~n20479;
  assign n20481 = n9331 & n12543;
  assign n20482 = n8418 & n12549;
  assign n20483 = n8860 & n12546;
  assign n20484 = ~n20482 & ~n20483;
  assign n20485 = ~n20481 & n20484;
  assign n20486 = n8421 & n15724;
  assign n20487 = n20485 & ~n20486;
  assign n20488 =  a[8]  & ~n20487;
  assign n20489 = ~n20487 & ~n20488;
  assign n20490 =  a[8]  & ~n20488;
  assign n20491 = ~n20489 & ~n20490;
  assign n20492 = ~n20046 & ~n20050;
  assign n20493 = ~n20049 & ~n20050;
  assign n20494 = ~n20492 & ~n20493;
  assign n20495 = ~n20491 & ~n20494;
  assign n20496 = ~n20491 & ~n20495;
  assign n20497 = ~n20494 & ~n20495;
  assign n20498 = ~n20496 & ~n20497;
  assign n20499 = n9331 & n12546;
  assign n20500 = n8418 & n12552;
  assign n20501 = n8860 & n12549;
  assign n20502 = ~n20500 & ~n20501;
  assign n20503 = ~n20499 & n20502;
  assign n20504 = n8421 & ~n15356;
  assign n20505 = n20503 & ~n20504;
  assign n20506 =  a[8]  & ~n20505;
  assign n20507 = ~n20505 & ~n20506;
  assign n20508 =  a[8]  & ~n20506;
  assign n20509 = ~n20507 & ~n20508;
  assign n20510 = ~n20041 & ~n20045;
  assign n20511 = ~n20044 & ~n20045;
  assign n20512 = ~n20510 & ~n20511;
  assign n20513 = ~n20509 & ~n20512;
  assign n20514 = ~n20509 & ~n20513;
  assign n20515 = ~n20512 & ~n20513;
  assign n20516 = ~n20514 & ~n20515;
  assign n20517 = n19942 & n20039;
  assign n20518 = ~n20040 & ~n20517;
  assign n20519 = n9331 & n12549;
  assign n20520 = n8418 & n12555;
  assign n20521 = n8860 & n12552;
  assign n20522 = ~n20520 & ~n20521;
  assign n20523 = ~n20519 & n20522;
  assign n20524 = ~n8421 & n20523;
  assign n20525 = ~n15764 & n20523;
  assign n20526 = ~n20524 & ~n20525;
  assign n20527 =  a[8]  & ~n20526;
  assign n20528 = ~ a[8]  & n20526;
  assign n20529 = ~n20527 & ~n20528;
  assign n20530 = n20518 & ~n20529;
  assign n20531 = n20035 & ~n20037;
  assign n20532 = ~n20038 & ~n20531;
  assign n20533 = n9331 & n12552;
  assign n20534 = n8418 & n12558;
  assign n20535 = n8860 & n12555;
  assign n20536 = ~n20534 & ~n20535;
  assign n20537 = ~n20533 & n20536;
  assign n20538 = ~n8421 & n20537;
  assign n20539 = n15791 & n20537;
  assign n20540 = ~n20538 & ~n20539;
  assign n20541 =  a[8]  & ~n20540;
  assign n20542 = ~ a[8]  & n20540;
  assign n20543 = ~n20541 & ~n20542;
  assign n20544 = n20532 & ~n20543;
  assign n20545 = n19974 & n20033;
  assign n20546 = ~n20034 & ~n20545;
  assign n20547 = n9331 & n12555;
  assign n20548 = n8418 & n12561;
  assign n20549 = n8860 & n12558;
  assign n20550 = ~n20548 & ~n20549;
  assign n20551 = ~n20547 & n20550;
  assign n20552 = ~n8421 & n20551;
  assign n20553 = n15816 & n20551;
  assign n20554 = ~n20552 & ~n20553;
  assign n20555 =  a[8]  & ~n20554;
  assign n20556 = ~ a[8]  & n20554;
  assign n20557 = ~n20555 & ~n20556;
  assign n20558 = n20546 & ~n20557;
  assign n20559 = n9331 & n12558;
  assign n20560 = n8418 & n12564;
  assign n20561 = n8860 & n12561;
  assign n20562 = ~n20560 & ~n20561;
  assign n20563 = ~n20559 & n20562;
  assign n20564 = n8421 & n15847;
  assign n20565 = n20563 & ~n20564;
  assign n20566 =  a[8]  & ~n20565;
  assign n20567 = ~n20565 & ~n20566;
  assign n20568 =  a[8]  & ~n20566;
  assign n20569 = ~n20567 & ~n20568;
  assign n20570 = n20029 & ~n20031;
  assign n20571 = ~n20032 & ~n20570;
  assign n20572 = ~n20569 & n20571;
  assign n20573 = ~n20569 & ~n20572;
  assign n20574 = n20571 & ~n20572;
  assign n20575 = ~n20573 & ~n20574;
  assign n20576 = ~n20016 & ~n20028;
  assign n20577 = ~n20027 & ~n20028;
  assign n20578 = ~n20576 & ~n20577;
  assign n20579 = n9331 & n12561;
  assign n20580 = n8418 & n12567;
  assign n20581 = n8860 & n12564;
  assign n20582 = ~n20580 & ~n20581;
  assign n20583 = ~n20579 & n20582;
  assign n20584 = ~n8421 & n20583;
  assign n20585 = n15905 & n20583;
  assign n20586 = ~n20584 & ~n20585;
  assign n20587 =  a[8]  & ~n20586;
  assign n20588 = ~ a[8]  & n20586;
  assign n20589 = ~n20587 & ~n20588;
  assign n20590 = ~n20578 & ~n20589;
  assign n20591 = n9331 & n12564;
  assign n20592 = n8418 & n12571;
  assign n20593 = n8860 & n12567;
  assign n20594 = ~n20592 & ~n20593;
  assign n20595 = ~n20591 & n20594;
  assign n20596 = n8421 & ~n15944;
  assign n20597 = n20595 & ~n20596;
  assign n20598 =  a[8]  & ~n20597;
  assign n20599 = ~n20597 & ~n20598;
  assign n20600 =  a[8]  & ~n20598;
  assign n20601 = ~n20599 & ~n20600;
  assign n20602 = ~n20000 & n20011;
  assign n20603 = ~n20012 & ~n20602;
  assign n20604 = ~n20601 & n20603;
  assign n20605 = ~n20601 & ~n20604;
  assign n20606 = n20603 & ~n20604;
  assign n20607 = ~n20605 & ~n20606;
  assign n20608 = n19997 & ~n19999;
  assign n20609 = ~n20000 & ~n20608;
  assign n20610 = n9331 & n12567;
  assign n20611 = n8418 & n12574;
  assign n20612 = n8860 & n12571;
  assign n20613 = ~n20611 & ~n20612;
  assign n20614 = ~n20610 & n20613;
  assign n20615 = ~n8421 & n20614;
  assign n20616 = ~n15989 & n20614;
  assign n20617 = ~n20615 & ~n20616;
  assign n20618 =  a[8]  & ~n20617;
  assign n20619 = ~ a[8]  & n20617;
  assign n20620 = ~n20618 & ~n20619;
  assign n20621 = n20609 & ~n20620;
  assign n20622 = n8860 & ~n12581;
  assign n20623 = n9331 & n12577;
  assign n20624 = ~n20622 & ~n20623;
  assign n20625 = n8421 & ~n16085;
  assign n20626 = n20624 & ~n20625;
  assign n20627 =  a[8]  & ~n20626;
  assign n20628 =  a[8]  & ~n20627;
  assign n20629 = ~n20626 & ~n20627;
  assign n20630 = ~n20628 & ~n20629;
  assign n20631 = ~n8416 & ~n12581;
  assign n20632 =  a[8]  & ~n20631;
  assign n20633 = ~n20630 & n20632;
  assign n20634 = n9331 & n12574;
  assign n20635 = n8418 & ~n12581;
  assign n20636 = n8860 & n12577;
  assign n20637 = ~n20635 & ~n20636;
  assign n20638 = ~n20634 & n20637;
  assign n20639 = ~n8421 & n20638;
  assign n20640 = n16094 & n20638;
  assign n20641 = ~n20639 & ~n20640;
  assign n20642 =  a[8]  & ~n20641;
  assign n20643 = ~ a[8]  & n20641;
  assign n20644 = ~n20642 & ~n20643;
  assign n20645 = n20633 & ~n20644;
  assign n20646 = n19998 & n20645;
  assign n20647 = n20645 & ~n20646;
  assign n20648 = n19998 & ~n20646;
  assign n20649 = ~n20647 & ~n20648;
  assign n20650 = n9331 & n12571;
  assign n20651 = n8418 & n12577;
  assign n20652 = n8860 & n12574;
  assign n20653 = ~n20651 & ~n20652;
  assign n20654 = ~n20650 & n20653;
  assign n20655 = n8421 & n16013;
  assign n20656 = n20654 & ~n20655;
  assign n20657 =  a[8]  & ~n20656;
  assign n20658 =  a[8]  & ~n20657;
  assign n20659 = ~n20656 & ~n20657;
  assign n20660 = ~n20658 & ~n20659;
  assign n20661 = ~n20649 & ~n20660;
  assign n20662 = ~n20646 & ~n20661;
  assign n20663 = ~n20609 & n20620;
  assign n20664 = ~n20621 & ~n20663;
  assign n20665 = ~n20662 & n20664;
  assign n20666 = ~n20621 & ~n20665;
  assign n20667 = ~n20607 & ~n20666;
  assign n20668 = ~n20604 & ~n20667;
  assign n20669 = n20578 & n20589;
  assign n20670 = ~n20590 & ~n20669;
  assign n20671 = ~n20668 & n20670;
  assign n20672 = ~n20590 & ~n20671;
  assign n20673 = ~n20575 & ~n20672;
  assign n20674 = ~n20572 & ~n20673;
  assign n20675 = n20546 & ~n20558;
  assign n20676 = ~n20557 & ~n20558;
  assign n20677 = ~n20675 & ~n20676;
  assign n20678 = ~n20674 & ~n20677;
  assign n20679 = ~n20558 & ~n20678;
  assign n20680 = n20532 & ~n20544;
  assign n20681 = ~n20543 & ~n20544;
  assign n20682 = ~n20680 & ~n20681;
  assign n20683 = ~n20679 & ~n20682;
  assign n20684 = ~n20544 & ~n20683;
  assign n20685 = ~n20518 & n20529;
  assign n20686 = ~n20530 & ~n20685;
  assign n20687 = ~n20684 & n20686;
  assign n20688 = ~n20530 & ~n20687;
  assign n20689 = ~n20516 & ~n20688;
  assign n20690 = ~n20513 & ~n20689;
  assign n20691 = ~n20498 & ~n20690;
  assign n20692 = ~n20495 & ~n20691;
  assign n20693 = ~n20480 & ~n20692;
  assign n20694 = ~n20477 & ~n20693;
  assign n20695 = n20451 & ~n20463;
  assign n20696 = ~n20462 & ~n20463;
  assign n20697 = ~n20695 & ~n20696;
  assign n20698 = ~n20694 & ~n20697;
  assign n20699 = ~n20463 & ~n20698;
  assign n20700 = n20437 & ~n20449;
  assign n20701 = ~n20448 & ~n20449;
  assign n20702 = ~n20700 & ~n20701;
  assign n20703 = ~n20699 & ~n20702;
  assign n20704 = ~n20449 & ~n20703;
  assign n20705 = ~n20423 & n20434;
  assign n20706 = ~n20435 & ~n20705;
  assign n20707 = ~n20704 & n20706;
  assign n20708 = ~n20435 & ~n20707;
  assign n20709 = ~n20421 & ~n20708;
  assign n20710 = ~n20418 & ~n20709;
  assign n20711 = ~n20403 & ~n20710;
  assign n20712 = ~n20400 & ~n20711;
  assign n20713 = ~n20385 & ~n20712;
  assign n20714 = ~n20382 & ~n20713;
  assign n20715 = n20356 & ~n20368;
  assign n20716 = ~n20367 & ~n20368;
  assign n20717 = ~n20715 & ~n20716;
  assign n20718 = ~n20714 & ~n20717;
  assign n20719 = ~n20368 & ~n20718;
  assign n20720 = n20342 & ~n20354;
  assign n20721 = ~n20353 & ~n20354;
  assign n20722 = ~n20720 & ~n20721;
  assign n20723 = ~n20719 & ~n20722;
  assign n20724 = ~n20354 & ~n20723;
  assign n20725 = ~n20328 & n20339;
  assign n20726 = ~n20340 & ~n20725;
  assign n20727 = ~n20724 & n20726;
  assign n20728 = ~n20340 & ~n20727;
  assign n20729 = ~n20326 & ~n20728;
  assign n20730 = ~n20323 & ~n20729;
  assign n20731 = ~n20308 & ~n20730;
  assign n20732 = ~n20305 & ~n20731;
  assign n20733 = n20279 & ~n20291;
  assign n20734 = ~n20290 & ~n20291;
  assign n20735 = ~n20733 & ~n20734;
  assign n20736 = ~n20732 & ~n20735;
  assign n20737 = ~n20291 & ~n20736;
  assign n20738 = n20265 & ~n20277;
  assign n20739 = ~n20276 & ~n20277;
  assign n20740 = ~n20738 & ~n20739;
  assign n20741 = ~n20737 & ~n20740;
  assign n20742 = ~n20277 & ~n20741;
  assign n20743 = n20251 & ~n20263;
  assign n20744 = ~n20262 & ~n20263;
  assign n20745 = ~n20743 & ~n20744;
  assign n20746 = ~n20742 & ~n20745;
  assign n20747 = ~n20263 & ~n20746;
  assign n20748 = n20237 & ~n20249;
  assign n20749 = ~n20248 & ~n20249;
  assign n20750 = ~n20748 & ~n20749;
  assign n20751 = ~n20747 & ~n20750;
  assign n20752 = ~n20249 & ~n20751;
  assign n20753 = n20223 & ~n20235;
  assign n20754 = ~n20234 & ~n20235;
  assign n20755 = ~n20753 & ~n20754;
  assign n20756 = ~n20752 & ~n20755;
  assign n20757 = ~n20235 & ~n20756;
  assign n20758 = n20209 & ~n20221;
  assign n20759 = ~n20220 & ~n20221;
  assign n20760 = ~n20758 & ~n20759;
  assign n20761 = ~n20757 & ~n20760;
  assign n20762 = ~n20221 & ~n20761;
  assign n20763 = n20195 & ~n20207;
  assign n20764 = ~n20206 & ~n20207;
  assign n20765 = ~n20763 & ~n20764;
  assign n20766 = ~n20762 & ~n20765;
  assign n20767 = ~n20207 & ~n20766;
  assign n20768 = n20181 & ~n20193;
  assign n20769 = ~n20192 & ~n20193;
  assign n20770 = ~n20768 & ~n20769;
  assign n20771 = ~n20767 & ~n20770;
  assign n20772 = ~n20193 & ~n20771;
  assign n20773 = n20167 & ~n20179;
  assign n20774 = ~n20178 & ~n20179;
  assign n20775 = ~n20773 & ~n20774;
  assign n20776 = ~n20772 & ~n20775;
  assign n20777 = ~n20179 & ~n20776;
  assign n20778 = ~n20153 & n20164;
  assign n20779 = ~n20165 & ~n20778;
  assign n20780 = ~n20777 & n20779;
  assign n20781 = ~n20165 & ~n20780;
  assign n20782 = ~n20151 & ~n20781;
  assign n20783 = n20151 & n20781;
  assign n20784 = ~n20782 & ~n20783;
  assign n20785 = n71 & n13941;
  assign n20786 = n9867 & n13633;
  assign n20787 = n10434 & ~n13627;
  assign n20788 = ~n20786 & ~n20787;
  assign n20789 = ~n20785 & n20788;
  assign n20790 = n9870 & n14136;
  assign n20791 = n20789 & ~n20790;
  assign n20792 =  a[5]  & ~n20791;
  assign n20793 =  a[5]  & ~n20792;
  assign n20794 = ~n20791 & ~n20792;
  assign n20795 = ~n20793 & ~n20794;
  assign n20796 = n20784 & ~n20795;
  assign n20797 = ~n20782 & ~n20796;
  assign n20798 = ~n20148 & ~n20797;
  assign n20799 = n20148 & n20797;
  assign n20800 = ~n20798 & ~n20799;
  assign n20801 = n20784 & ~n20796;
  assign n20802 = ~n20795 & ~n20796;
  assign n20803 = ~n20801 & ~n20802;
  assign n20804 = n71 & ~n13627;
  assign n20805 = n9867 & n13630;
  assign n20806 = n10434 & n13633;
  assign n20807 = ~n20805 & ~n20806;
  assign n20808 = ~n20804 & n20807;
  assign n20809 = n9870 & ~n13654;
  assign n20810 = n20808 & ~n20809;
  assign n20811 =  a[5]  & ~n20810;
  assign n20812 = ~n20810 & ~n20811;
  assign n20813 =  a[5]  & ~n20811;
  assign n20814 = ~n20812 & ~n20813;
  assign n20815 = n20777 & ~n20779;
  assign n20816 = ~n20780 & ~n20815;
  assign n20817 = ~n20814 & n20816;
  assign n20818 = ~n20814 & ~n20817;
  assign n20819 = n20816 & ~n20817;
  assign n20820 = ~n20818 & ~n20819;
  assign n20821 = ~n11715 & ~n11727;
  assign n20822 = ~n13438 & ~n20821;
  assign n20823 = n11055 & n13941;
  assign n20824 = ~n20822 & ~n20823;
  assign n20825 = n11057 & ~n13951;
  assign n20826 = n20824 & ~n20825;
  assign n20827 =  a[2]  & ~n20826;
  assign n20828 =  a[2]  & ~n20827;
  assign n20829 = ~n20826 & ~n20827;
  assign n20830 = ~n20828 & ~n20829;
  assign n20831 = ~n20820 & ~n20830;
  assign n20832 = ~n20817 & ~n20831;
  assign n20833 = ~n20803 & ~n20832;
  assign n20834 = n20803 & n20832;
  assign n20835 = ~n20833 & ~n20834;
  assign n20836 = ~n20820 & ~n20831;
  assign n20837 = ~n20830 & ~n20831;
  assign n20838 = ~n20836 & ~n20837;
  assign n20839 = n71 & n13633;
  assign n20840 = n9867 & n13597;
  assign n20841 = n10434 & n13630;
  assign n20842 = ~n20840 & ~n20841;
  assign n20843 = ~n20839 & n20842;
  assign n20844 = n9870 & n13929;
  assign n20845 = n20843 & ~n20844;
  assign n20846 =  a[5]  & ~n20845;
  assign n20847 = ~n20845 & ~n20846;
  assign n20848 =  a[5]  & ~n20846;
  assign n20849 = ~n20847 & ~n20848;
  assign n20850 = ~n20772 & ~n20776;
  assign n20851 = ~n20775 & ~n20776;
  assign n20852 = ~n20850 & ~n20851;
  assign n20853 = ~n20849 & ~n20852;
  assign n20854 = ~n20849 & ~n20853;
  assign n20855 = ~n20852 & ~n20853;
  assign n20856 = ~n20854 & ~n20855;
  assign n20857 = n71 & n13630;
  assign n20858 = n9867 & n13515;
  assign n20859 = n10434 & n13597;
  assign n20860 = ~n20858 & ~n20859;
  assign n20861 = ~n20857 & n20860;
  assign n20862 = n9870 & n13976;
  assign n20863 = n20861 & ~n20862;
  assign n20864 =  a[5]  & ~n20863;
  assign n20865 = ~n20863 & ~n20864;
  assign n20866 =  a[5]  & ~n20864;
  assign n20867 = ~n20865 & ~n20866;
  assign n20868 = ~n20767 & ~n20771;
  assign n20869 = ~n20770 & ~n20771;
  assign n20870 = ~n20868 & ~n20869;
  assign n20871 = ~n20867 & ~n20870;
  assign n20872 = ~n20867 & ~n20871;
  assign n20873 = ~n20870 & ~n20871;
  assign n20874 = ~n20872 & ~n20873;
  assign n20875 = n71 & n13597;
  assign n20876 = n9867 & n13521;
  assign n20877 = n10434 & n13515;
  assign n20878 = ~n20876 & ~n20877;
  assign n20879 = ~n20875 & n20878;
  assign n20880 = n9870 & ~n13612;
  assign n20881 = n20879 & ~n20880;
  assign n20882 =  a[5]  & ~n20881;
  assign n20883 = ~n20881 & ~n20882;
  assign n20884 =  a[5]  & ~n20882;
  assign n20885 = ~n20883 & ~n20884;
  assign n20886 = ~n20762 & ~n20766;
  assign n20887 = ~n20765 & ~n20766;
  assign n20888 = ~n20886 & ~n20887;
  assign n20889 = ~n20885 & ~n20888;
  assign n20890 = ~n20885 & ~n20889;
  assign n20891 = ~n20888 & ~n20889;
  assign n20892 = ~n20890 & ~n20891;
  assign n20893 = n71 & n13515;
  assign n20894 = n9867 & n13518;
  assign n20895 = n10434 & n13521;
  assign n20896 = ~n20894 & ~n20895;
  assign n20897 = ~n20893 & n20896;
  assign n20898 = n9870 & n13541;
  assign n20899 = n20897 & ~n20898;
  assign n20900 =  a[5]  & ~n20899;
  assign n20901 = ~n20899 & ~n20900;
  assign n20902 =  a[5]  & ~n20900;
  assign n20903 = ~n20901 & ~n20902;
  assign n20904 = ~n20757 & ~n20761;
  assign n20905 = ~n20760 & ~n20761;
  assign n20906 = ~n20904 & ~n20905;
  assign n20907 = ~n20903 & ~n20906;
  assign n20908 = ~n20903 & ~n20907;
  assign n20909 = ~n20906 & ~n20907;
  assign n20910 = ~n20908 & ~n20909;
  assign n20911 = n71 & n13521;
  assign n20912 = n9867 & n13491;
  assign n20913 = n10434 & n13518;
  assign n20914 = ~n20912 & ~n20913;
  assign n20915 = ~n20911 & n20914;
  assign n20916 = n9870 & ~n13909;
  assign n20917 = n20915 & ~n20916;
  assign n20918 =  a[5]  & ~n20917;
  assign n20919 = ~n20917 & ~n20918;
  assign n20920 =  a[5]  & ~n20918;
  assign n20921 = ~n20919 & ~n20920;
  assign n20922 = ~n20752 & ~n20756;
  assign n20923 = ~n20755 & ~n20756;
  assign n20924 = ~n20922 & ~n20923;
  assign n20925 = ~n20921 & ~n20924;
  assign n20926 = ~n20921 & ~n20925;
  assign n20927 = ~n20924 & ~n20925;
  assign n20928 = ~n20926 & ~n20927;
  assign n20929 = n71 & n13518;
  assign n20930 = n9867 & n12889;
  assign n20931 = n10434 & n13491;
  assign n20932 = ~n20930 & ~n20931;
  assign n20933 = ~n20929 & n20932;
  assign n20934 = n9870 & n13584;
  assign n20935 = n20933 & ~n20934;
  assign n20936 =  a[5]  & ~n20935;
  assign n20937 = ~n20935 & ~n20936;
  assign n20938 =  a[5]  & ~n20936;
  assign n20939 = ~n20937 & ~n20938;
  assign n20940 = ~n20747 & ~n20751;
  assign n20941 = ~n20750 & ~n20751;
  assign n20942 = ~n20940 & ~n20941;
  assign n20943 = ~n20939 & ~n20942;
  assign n20944 = ~n20939 & ~n20943;
  assign n20945 = ~n20942 & ~n20943;
  assign n20946 = ~n20944 & ~n20945;
  assign n20947 = n71 & n13491;
  assign n20948 = n9867 & n12769;
  assign n20949 = n10434 & n12889;
  assign n20950 = ~n20948 & ~n20949;
  assign n20951 = ~n20947 & n20950;
  assign n20952 = n9870 & ~n13503;
  assign n20953 = n20951 & ~n20952;
  assign n20954 =  a[5]  & ~n20953;
  assign n20955 = ~n20953 & ~n20954;
  assign n20956 =  a[5]  & ~n20954;
  assign n20957 = ~n20955 & ~n20956;
  assign n20958 = ~n20742 & ~n20746;
  assign n20959 = ~n20745 & ~n20746;
  assign n20960 = ~n20958 & ~n20959;
  assign n20961 = ~n20957 & ~n20960;
  assign n20962 = ~n20957 & ~n20961;
  assign n20963 = ~n20960 & ~n20961;
  assign n20964 = ~n20962 & ~n20963;
  assign n20965 = n71 & n12889;
  assign n20966 = n9867 & n12502;
  assign n20967 = n10434 & n12769;
  assign n20968 = ~n20966 & ~n20967;
  assign n20969 = ~n20965 & n20968;
  assign n20970 = n9870 & n12895;
  assign n20971 = n20969 & ~n20970;
  assign n20972 =  a[5]  & ~n20971;
  assign n20973 = ~n20971 & ~n20972;
  assign n20974 =  a[5]  & ~n20972;
  assign n20975 = ~n20973 & ~n20974;
  assign n20976 = ~n20737 & ~n20741;
  assign n20977 = ~n20740 & ~n20741;
  assign n20978 = ~n20976 & ~n20977;
  assign n20979 = ~n20975 & ~n20978;
  assign n20980 = ~n20975 & ~n20979;
  assign n20981 = ~n20978 & ~n20979;
  assign n20982 = ~n20980 & ~n20981;
  assign n20983 = n71 & n12769;
  assign n20984 = n9867 & n12370;
  assign n20985 = n10434 & n12502;
  assign n20986 = ~n20984 & ~n20985;
  assign n20987 = ~n20983 & n20986;
  assign n20988 = n9870 & n12999;
  assign n20989 = n20987 & ~n20988;
  assign n20990 =  a[5]  & ~n20989;
  assign n20991 = ~n20989 & ~n20990;
  assign n20992 =  a[5]  & ~n20990;
  assign n20993 = ~n20991 & ~n20992;
  assign n20994 = ~n20732 & ~n20736;
  assign n20995 = ~n20735 & ~n20736;
  assign n20996 = ~n20994 & ~n20995;
  assign n20997 = ~n20993 & ~n20996;
  assign n20998 = ~n20993 & ~n20997;
  assign n20999 = ~n20996 & ~n20997;
  assign n21000 = ~n20998 & ~n20999;
  assign n21001 = n20308 & n20730;
  assign n21002 = ~n20731 & ~n21001;
  assign n21003 = n71 & n12502;
  assign n21004 = n9867 & n12505;
  assign n21005 = n10434 & n12370;
  assign n21006 = ~n21004 & ~n21005;
  assign n21007 = ~n21003 & n21006;
  assign n21008 = ~n9870 & n21007;
  assign n21009 = n13736 & n21007;
  assign n21010 = ~n21008 & ~n21009;
  assign n21011 =  a[5]  & ~n21010;
  assign n21012 = ~ a[5]  & n21010;
  assign n21013 = ~n21011 & ~n21012;
  assign n21014 = n21002 & ~n21013;
  assign n21015 = n20326 & n20728;
  assign n21016 = ~n20729 & ~n21015;
  assign n21017 = n71 & n12370;
  assign n21018 = n9867 & n12508;
  assign n21019 = n10434 & n12505;
  assign n21020 = ~n21018 & ~n21019;
  assign n21021 = ~n21017 & n21020;
  assign n21022 = ~n9870 & n21021;
  assign n21023 = n13748 & n21021;
  assign n21024 = ~n21022 & ~n21023;
  assign n21025 =  a[5]  & ~n21024;
  assign n21026 = ~ a[5]  & n21024;
  assign n21027 = ~n21025 & ~n21026;
  assign n21028 = n21016 & ~n21027;
  assign n21029 = n71 & n12505;
  assign n21030 = n9867 & n12513;
  assign n21031 = n10434 & n12508;
  assign n21032 = ~n21030 & ~n21031;
  assign n21033 = ~n21029 & n21032;
  assign n21034 = n9870 & ~n14051;
  assign n21035 = n21033 & ~n21034;
  assign n21036 =  a[5]  & ~n21035;
  assign n21037 = ~n21035 & ~n21036;
  assign n21038 =  a[5]  & ~n21036;
  assign n21039 = ~n21037 & ~n21038;
  assign n21040 = n20724 & ~n20726;
  assign n21041 = ~n20727 & ~n21040;
  assign n21042 = ~n21039 & n21041;
  assign n21043 = ~n21039 & ~n21042;
  assign n21044 = n21041 & ~n21042;
  assign n21045 = ~n21043 & ~n21044;
  assign n21046 = n71 & n12508;
  assign n21047 = n9867 & n12511;
  assign n21048 = n10434 & n12513;
  assign n21049 = ~n21047 & ~n21048;
  assign n21050 = ~n21046 & n21049;
  assign n21051 = n9870 & n13863;
  assign n21052 = n21050 & ~n21051;
  assign n21053 =  a[5]  & ~n21052;
  assign n21054 = ~n21052 & ~n21053;
  assign n21055 =  a[5]  & ~n21053;
  assign n21056 = ~n21054 & ~n21055;
  assign n21057 = ~n20719 & ~n20723;
  assign n21058 = ~n20722 & ~n20723;
  assign n21059 = ~n21057 & ~n21058;
  assign n21060 = ~n21056 & ~n21059;
  assign n21061 = ~n21056 & ~n21060;
  assign n21062 = ~n21059 & ~n21060;
  assign n21063 = ~n21061 & ~n21062;
  assign n21064 = n71 & n12513;
  assign n21065 = n9867 & n12516;
  assign n21066 = n10434 & n12511;
  assign n21067 = ~n21065 & ~n21066;
  assign n21068 = ~n21064 & n21067;
  assign n21069 = n9870 & n14177;
  assign n21070 = n21068 & ~n21069;
  assign n21071 =  a[5]  & ~n21070;
  assign n21072 = ~n21070 & ~n21071;
  assign n21073 =  a[5]  & ~n21071;
  assign n21074 = ~n21072 & ~n21073;
  assign n21075 = ~n20714 & ~n20718;
  assign n21076 = ~n20717 & ~n20718;
  assign n21077 = ~n21075 & ~n21076;
  assign n21078 = ~n21074 & ~n21077;
  assign n21079 = ~n21074 & ~n21078;
  assign n21080 = ~n21077 & ~n21078;
  assign n21081 = ~n21079 & ~n21080;
  assign n21082 = n20385 & n20712;
  assign n21083 = ~n20713 & ~n21082;
  assign n21084 = n71 & n12511;
  assign n21085 = n9867 & n12519;
  assign n21086 = n10434 & n12516;
  assign n21087 = ~n21085 & ~n21086;
  assign n21088 = ~n21084 & n21087;
  assign n21089 = ~n9870 & n21088;
  assign n21090 = n14233 & n21088;
  assign n21091 = ~n21089 & ~n21090;
  assign n21092 =  a[5]  & ~n21091;
  assign n21093 = ~ a[5]  & n21091;
  assign n21094 = ~n21092 & ~n21093;
  assign n21095 = n21083 & ~n21094;
  assign n21096 = n20403 & n20710;
  assign n21097 = ~n20711 & ~n21096;
  assign n21098 = n71 & n12516;
  assign n21099 = n9867 & n12522;
  assign n21100 = n10434 & n12519;
  assign n21101 = ~n21099 & ~n21100;
  assign n21102 = ~n21098 & n21101;
  assign n21103 = ~n9870 & n21102;
  assign n21104 = n14443 & n21102;
  assign n21105 = ~n21103 & ~n21104;
  assign n21106 =  a[5]  & ~n21105;
  assign n21107 = ~ a[5]  & n21105;
  assign n21108 = ~n21106 & ~n21107;
  assign n21109 = n21097 & ~n21108;
  assign n21110 = n20421 & n20708;
  assign n21111 = ~n20709 & ~n21110;
  assign n21112 = n71 & n12519;
  assign n21113 = n9867 & n12525;
  assign n21114 = n10434 & n12522;
  assign n21115 = ~n21113 & ~n21114;
  assign n21116 = ~n21112 & n21115;
  assign n21117 = ~n9870 & n21116;
  assign n21118 = ~n14454 & n21116;
  assign n21119 = ~n21117 & ~n21118;
  assign n21120 =  a[5]  & ~n21119;
  assign n21121 = ~ a[5]  & n21119;
  assign n21122 = ~n21120 & ~n21121;
  assign n21123 = n21111 & ~n21122;
  assign n21124 = n71 & n12522;
  assign n21125 = n9867 & n12528;
  assign n21126 = n10434 & n12525;
  assign n21127 = ~n21125 & ~n21126;
  assign n21128 = ~n21124 & n21127;
  assign n21129 = n9870 & n14837;
  assign n21130 = n21128 & ~n21129;
  assign n21131 =  a[5]  & ~n21130;
  assign n21132 = ~n21130 & ~n21131;
  assign n21133 =  a[5]  & ~n21131;
  assign n21134 = ~n21132 & ~n21133;
  assign n21135 = n20704 & ~n20706;
  assign n21136 = ~n20707 & ~n21135;
  assign n21137 = ~n21134 & n21136;
  assign n21138 = ~n21134 & ~n21137;
  assign n21139 = n21136 & ~n21137;
  assign n21140 = ~n21138 & ~n21139;
  assign n21141 = n71 & n12525;
  assign n21142 = n9867 & n12531;
  assign n21143 = n10434 & n12528;
  assign n21144 = ~n21142 & ~n21143;
  assign n21145 = ~n21141 & n21144;
  assign n21146 = n9870 & n14608;
  assign n21147 = n21145 & ~n21146;
  assign n21148 =  a[5]  & ~n21147;
  assign n21149 = ~n21147 & ~n21148;
  assign n21150 =  a[5]  & ~n21148;
  assign n21151 = ~n21149 & ~n21150;
  assign n21152 = ~n20699 & ~n20703;
  assign n21153 = ~n20702 & ~n20703;
  assign n21154 = ~n21152 & ~n21153;
  assign n21155 = ~n21151 & ~n21154;
  assign n21156 = ~n21151 & ~n21155;
  assign n21157 = ~n21154 & ~n21155;
  assign n21158 = ~n21156 & ~n21157;
  assign n21159 = n71 & n12528;
  assign n21160 = n9867 & n12534;
  assign n21161 = n10434 & n12531;
  assign n21162 = ~n21160 & ~n21161;
  assign n21163 = ~n21159 & n21162;
  assign n21164 = n9870 & ~n15003;
  assign n21165 = n21163 & ~n21164;
  assign n21166 =  a[5]  & ~n21165;
  assign n21167 = ~n21165 & ~n21166;
  assign n21168 =  a[5]  & ~n21166;
  assign n21169 = ~n21167 & ~n21168;
  assign n21170 = ~n20694 & ~n20698;
  assign n21171 = ~n20697 & ~n20698;
  assign n21172 = ~n21170 & ~n21171;
  assign n21173 = ~n21169 & ~n21172;
  assign n21174 = ~n21169 & ~n21173;
  assign n21175 = ~n21172 & ~n21173;
  assign n21176 = ~n21174 & ~n21175;
  assign n21177 = n20480 & n20692;
  assign n21178 = ~n20693 & ~n21177;
  assign n21179 = n71 & n12531;
  assign n21180 = n9867 & n12537;
  assign n21181 = n10434 & n12534;
  assign n21182 = ~n21180 & ~n21181;
  assign n21183 = ~n21179 & n21182;
  assign n21184 = ~n9870 & n21183;
  assign n21185 = ~n15255 & n21183;
  assign n21186 = ~n21184 & ~n21185;
  assign n21187 =  a[5]  & ~n21186;
  assign n21188 = ~ a[5]  & n21186;
  assign n21189 = ~n21187 & ~n21188;
  assign n21190 = n21178 & ~n21189;
  assign n21191 = n20498 & n20690;
  assign n21192 = ~n20691 & ~n21191;
  assign n21193 = n71 & n12534;
  assign n21194 = n9867 & n12540;
  assign n21195 = n10434 & n12537;
  assign n21196 = ~n21194 & ~n21195;
  assign n21197 = ~n21193 & n21196;
  assign n21198 = ~n9870 & n21197;
  assign n21199 = n15096 & n21197;
  assign n21200 = ~n21198 & ~n21199;
  assign n21201 =  a[5]  & ~n21200;
  assign n21202 = ~ a[5]  & n21200;
  assign n21203 = ~n21201 & ~n21202;
  assign n21204 = n21192 & ~n21203;
  assign n21205 = n20516 & n20688;
  assign n21206 = ~n20689 & ~n21205;
  assign n21207 = n71 & n12537;
  assign n21208 = n9867 & n12543;
  assign n21209 = n10434 & n12540;
  assign n21210 = ~n21208 & ~n21209;
  assign n21211 = ~n21207 & n21210;
  assign n21212 = ~n9870 & n21211;
  assign n21213 = n15385 & n21211;
  assign n21214 = ~n21212 & ~n21213;
  assign n21215 =  a[5]  & ~n21214;
  assign n21216 = ~ a[5]  & n21214;
  assign n21217 = ~n21215 & ~n21216;
  assign n21218 = n21206 & ~n21217;
  assign n21219 = n71 & n12540;
  assign n21220 = n9867 & n12546;
  assign n21221 = n10434 & n12543;
  assign n21222 = ~n21220 & ~n21221;
  assign n21223 = ~n21219 & n21222;
  assign n21224 = n9870 & ~n15708;
  assign n21225 = n21223 & ~n21224;
  assign n21226 =  a[5]  & ~n21225;
  assign n21227 = ~n21225 & ~n21226;
  assign n21228 =  a[5]  & ~n21226;
  assign n21229 = ~n21227 & ~n21228;
  assign n21230 = n20684 & ~n20686;
  assign n21231 = ~n20687 & ~n21230;
  assign n21232 = ~n21229 & n21231;
  assign n21233 = ~n21229 & ~n21232;
  assign n21234 = n21231 & ~n21232;
  assign n21235 = ~n21233 & ~n21234;
  assign n21236 = n71 & n12543;
  assign n21237 = n9867 & n12549;
  assign n21238 = n10434 & n12546;
  assign n21239 = ~n21237 & ~n21238;
  assign n21240 = ~n21236 & n21239;
  assign n21241 = n9870 & n15724;
  assign n21242 = n21240 & ~n21241;
  assign n21243 =  a[5]  & ~n21242;
  assign n21244 = ~n21242 & ~n21243;
  assign n21245 =  a[5]  & ~n21243;
  assign n21246 = ~n21244 & ~n21245;
  assign n21247 = ~n20679 & ~n20683;
  assign n21248 = ~n20682 & ~n20683;
  assign n21249 = ~n21247 & ~n21248;
  assign n21250 = ~n21246 & ~n21249;
  assign n21251 = ~n21246 & ~n21250;
  assign n21252 = ~n21249 & ~n21250;
  assign n21253 = ~n21251 & ~n21252;
  assign n21254 = n71 & n12546;
  assign n21255 = n9867 & n12552;
  assign n21256 = n10434 & n12549;
  assign n21257 = ~n21255 & ~n21256;
  assign n21258 = ~n21254 & n21257;
  assign n21259 = n9870 & ~n15356;
  assign n21260 = n21258 & ~n21259;
  assign n21261 =  a[5]  & ~n21260;
  assign n21262 = ~n21260 & ~n21261;
  assign n21263 =  a[5]  & ~n21261;
  assign n21264 = ~n21262 & ~n21263;
  assign n21265 = ~n20674 & ~n20678;
  assign n21266 = ~n20677 & ~n20678;
  assign n21267 = ~n21265 & ~n21266;
  assign n21268 = ~n21264 & ~n21267;
  assign n21269 = ~n21264 & ~n21268;
  assign n21270 = ~n21267 & ~n21268;
  assign n21271 = ~n21269 & ~n21270;
  assign n21272 = n20575 & n20672;
  assign n21273 = ~n20673 & ~n21272;
  assign n21274 = n71 & n12549;
  assign n21275 = n9867 & n12555;
  assign n21276 = n10434 & n12552;
  assign n21277 = ~n21275 & ~n21276;
  assign n21278 = ~n21274 & n21277;
  assign n21279 = ~n9870 & n21278;
  assign n21280 = ~n15764 & n21278;
  assign n21281 = ~n21279 & ~n21280;
  assign n21282 =  a[5]  & ~n21281;
  assign n21283 = ~ a[5]  & n21281;
  assign n21284 = ~n21282 & ~n21283;
  assign n21285 = n21273 & ~n21284;
  assign n21286 = n20668 & ~n20670;
  assign n21287 = ~n20671 & ~n21286;
  assign n21288 = n71 & n12552;
  assign n21289 = n9867 & n12558;
  assign n21290 = n10434 & n12555;
  assign n21291 = ~n21289 & ~n21290;
  assign n21292 = ~n21288 & n21291;
  assign n21293 = ~n9870 & n21292;
  assign n21294 = n15791 & n21292;
  assign n21295 = ~n21293 & ~n21294;
  assign n21296 =  a[5]  & ~n21295;
  assign n21297 = ~ a[5]  & n21295;
  assign n21298 = ~n21296 & ~n21297;
  assign n21299 = n21287 & ~n21298;
  assign n21300 = n20607 & n20666;
  assign n21301 = ~n20667 & ~n21300;
  assign n21302 = n71 & n12555;
  assign n21303 = n9867 & n12561;
  assign n21304 = n10434 & n12558;
  assign n21305 = ~n21303 & ~n21304;
  assign n21306 = ~n21302 & n21305;
  assign n21307 = ~n9870 & n21306;
  assign n21308 = n15816 & n21306;
  assign n21309 = ~n21307 & ~n21308;
  assign n21310 =  a[5]  & ~n21309;
  assign n21311 = ~ a[5]  & n21309;
  assign n21312 = ~n21310 & ~n21311;
  assign n21313 = n21301 & ~n21312;
  assign n21314 = n71 & n12558;
  assign n21315 = n9867 & n12564;
  assign n21316 = n10434 & n12561;
  assign n21317 = ~n21315 & ~n21316;
  assign n21318 = ~n21314 & n21317;
  assign n21319 = n9870 & n15847;
  assign n21320 = n21318 & ~n21319;
  assign n21321 =  a[5]  & ~n21320;
  assign n21322 = ~n21320 & ~n21321;
  assign n21323 =  a[5]  & ~n21321;
  assign n21324 = ~n21322 & ~n21323;
  assign n21325 = n20662 & ~n20664;
  assign n21326 = ~n20665 & ~n21325;
  assign n21327 = ~n21324 & n21326;
  assign n21328 = ~n21324 & ~n21327;
  assign n21329 = n21326 & ~n21327;
  assign n21330 = ~n21328 & ~n21329;
  assign n21331 = ~n20649 & ~n20661;
  assign n21332 = ~n20660 & ~n20661;
  assign n21333 = ~n21331 & ~n21332;
  assign n21334 = n71 & n12561;
  assign n21335 = n9867 & n12567;
  assign n21336 = n10434 & n12564;
  assign n21337 = ~n21335 & ~n21336;
  assign n21338 = ~n21334 & n21337;
  assign n21339 = ~n9870 & n21338;
  assign n21340 = n15905 & n21338;
  assign n21341 = ~n21339 & ~n21340;
  assign n21342 =  a[5]  & ~n21341;
  assign n21343 = ~ a[5]  & n21341;
  assign n21344 = ~n21342 & ~n21343;
  assign n21345 = ~n21333 & ~n21344;
  assign n21346 = n71 & n12564;
  assign n21347 = n9867 & n12571;
  assign n21348 = n10434 & n12567;
  assign n21349 = ~n21347 & ~n21348;
  assign n21350 = ~n21346 & n21349;
  assign n21351 = n9870 & ~n15944;
  assign n21352 = n21350 & ~n21351;
  assign n21353 =  a[5]  & ~n21352;
  assign n21354 = ~n21352 & ~n21353;
  assign n21355 =  a[5]  & ~n21353;
  assign n21356 = ~n21354 & ~n21355;
  assign n21357 = ~n20633 & n20644;
  assign n21358 = ~n20645 & ~n21357;
  assign n21359 = ~n21356 & n21358;
  assign n21360 = ~n21356 & ~n21359;
  assign n21361 = n21358 & ~n21359;
  assign n21362 = ~n21360 & ~n21361;
  assign n21363 = n20630 & ~n20632;
  assign n21364 = ~n20633 & ~n21363;
  assign n21365 = n71 & n12567;
  assign n21366 = n9867 & n12574;
  assign n21367 = n10434 & n12571;
  assign n21368 = ~n21366 & ~n21367;
  assign n21369 = ~n21365 & n21368;
  assign n21370 = ~n9870 & n21369;
  assign n21371 = ~n15989 & n21369;
  assign n21372 = ~n21370 & ~n21371;
  assign n21373 =  a[5]  & ~n21372;
  assign n21374 = ~ a[5]  & n21372;
  assign n21375 = ~n21373 & ~n21374;
  assign n21376 = n21364 & ~n21375;
  assign n21377 = n10434 & ~n12581;
  assign n21378 = n71 & n12577;
  assign n21379 = ~n21377 & ~n21378;
  assign n21380 = n9870 & ~n16085;
  assign n21381 = n21379 & ~n21380;
  assign n21382 =  a[5]  & ~n21381;
  assign n21383 =  a[5]  & ~n21382;
  assign n21384 = ~n21381 & ~n21382;
  assign n21385 = ~n21383 & ~n21384;
  assign n21386 = ~n70 & ~n12581;
  assign n21387 =  a[5]  & ~n21386;
  assign n21388 = ~n21385 & n21387;
  assign n21389 = n71 & n12574;
  assign n21390 = n9867 & ~n12581;
  assign n21391 = n10434 & n12577;
  assign n21392 = ~n21390 & ~n21391;
  assign n21393 = ~n21389 & n21392;
  assign n21394 = ~n9870 & n21393;
  assign n21395 = n16094 & n21393;
  assign n21396 = ~n21394 & ~n21395;
  assign n21397 =  a[5]  & ~n21396;
  assign n21398 = ~ a[5]  & n21396;
  assign n21399 = ~n21397 & ~n21398;
  assign n21400 = n21388 & ~n21399;
  assign n21401 = n20631 & n21400;
  assign n21402 = n21400 & ~n21401;
  assign n21403 = n20631 & ~n21401;
  assign n21404 = ~n21402 & ~n21403;
  assign n21405 = n71 & n12571;
  assign n21406 = n9867 & n12577;
  assign n21407 = n10434 & n12574;
  assign n21408 = ~n21406 & ~n21407;
  assign n21409 = ~n21405 & n21408;
  assign n21410 = n9870 & n16013;
  assign n21411 = n21409 & ~n21410;
  assign n21412 =  a[5]  & ~n21411;
  assign n21413 =  a[5]  & ~n21412;
  assign n21414 = ~n21411 & ~n21412;
  assign n21415 = ~n21413 & ~n21414;
  assign n21416 = ~n21404 & ~n21415;
  assign n21417 = ~n21401 & ~n21416;
  assign n21418 = ~n21364 & n21375;
  assign n21419 = ~n21376 & ~n21418;
  assign n21420 = ~n21417 & n21419;
  assign n21421 = ~n21376 & ~n21420;
  assign n21422 = ~n21362 & ~n21421;
  assign n21423 = ~n21359 & ~n21422;
  assign n21424 = n21333 & n21344;
  assign n21425 = ~n21345 & ~n21424;
  assign n21426 = ~n21423 & n21425;
  assign n21427 = ~n21345 & ~n21426;
  assign n21428 = ~n21330 & ~n21427;
  assign n21429 = ~n21327 & ~n21428;
  assign n21430 = n21301 & ~n21313;
  assign n21431 = ~n21312 & ~n21313;
  assign n21432 = ~n21430 & ~n21431;
  assign n21433 = ~n21429 & ~n21432;
  assign n21434 = ~n21313 & ~n21433;
  assign n21435 = n21287 & ~n21299;
  assign n21436 = ~n21298 & ~n21299;
  assign n21437 = ~n21435 & ~n21436;
  assign n21438 = ~n21434 & ~n21437;
  assign n21439 = ~n21299 & ~n21438;
  assign n21440 = ~n21273 & n21284;
  assign n21441 = ~n21285 & ~n21440;
  assign n21442 = ~n21439 & n21441;
  assign n21443 = ~n21285 & ~n21442;
  assign n21444 = ~n21271 & ~n21443;
  assign n21445 = ~n21268 & ~n21444;
  assign n21446 = ~n21253 & ~n21445;
  assign n21447 = ~n21250 & ~n21446;
  assign n21448 = ~n21235 & ~n21447;
  assign n21449 = ~n21232 & ~n21448;
  assign n21450 = n21206 & ~n21218;
  assign n21451 = ~n21217 & ~n21218;
  assign n21452 = ~n21450 & ~n21451;
  assign n21453 = ~n21449 & ~n21452;
  assign n21454 = ~n21218 & ~n21453;
  assign n21455 = n21192 & ~n21204;
  assign n21456 = ~n21203 & ~n21204;
  assign n21457 = ~n21455 & ~n21456;
  assign n21458 = ~n21454 & ~n21457;
  assign n21459 = ~n21204 & ~n21458;
  assign n21460 = ~n21178 & n21189;
  assign n21461 = ~n21190 & ~n21460;
  assign n21462 = ~n21459 & n21461;
  assign n21463 = ~n21190 & ~n21462;
  assign n21464 = ~n21176 & ~n21463;
  assign n21465 = ~n21173 & ~n21464;
  assign n21466 = ~n21158 & ~n21465;
  assign n21467 = ~n21155 & ~n21466;
  assign n21468 = ~n21140 & ~n21467;
  assign n21469 = ~n21137 & ~n21468;
  assign n21470 = n21111 & ~n21123;
  assign n21471 = ~n21122 & ~n21123;
  assign n21472 = ~n21470 & ~n21471;
  assign n21473 = ~n21469 & ~n21472;
  assign n21474 = ~n21123 & ~n21473;
  assign n21475 = n21097 & ~n21109;
  assign n21476 = ~n21108 & ~n21109;
  assign n21477 = ~n21475 & ~n21476;
  assign n21478 = ~n21474 & ~n21477;
  assign n21479 = ~n21109 & ~n21478;
  assign n21480 = ~n21083 & n21094;
  assign n21481 = ~n21095 & ~n21480;
  assign n21482 = ~n21479 & n21481;
  assign n21483 = ~n21095 & ~n21482;
  assign n21484 = ~n21081 & ~n21483;
  assign n21485 = ~n21078 & ~n21484;
  assign n21486 = ~n21063 & ~n21485;
  assign n21487 = ~n21060 & ~n21486;
  assign n21488 = ~n21045 & ~n21487;
  assign n21489 = ~n21042 & ~n21488;
  assign n21490 = n21016 & ~n21028;
  assign n21491 = ~n21027 & ~n21028;
  assign n21492 = ~n21490 & ~n21491;
  assign n21493 = ~n21489 & ~n21492;
  assign n21494 = ~n21028 & ~n21493;
  assign n21495 = ~n21002 & n21013;
  assign n21496 = ~n21014 & ~n21495;
  assign n21497 = ~n21494 & n21496;
  assign n21498 = ~n21014 & ~n21497;
  assign n21499 = ~n21000 & ~n21498;
  assign n21500 = ~n20997 & ~n21499;
  assign n21501 = ~n20982 & ~n21500;
  assign n21502 = ~n20979 & ~n21501;
  assign n21503 = ~n20964 & ~n21502;
  assign n21504 = ~n20961 & ~n21503;
  assign n21505 = ~n20946 & ~n21504;
  assign n21506 = ~n20943 & ~n21505;
  assign n21507 = ~n20928 & ~n21506;
  assign n21508 = ~n20925 & ~n21507;
  assign n21509 = ~n20910 & ~n21508;
  assign n21510 = ~n20907 & ~n21509;
  assign n21511 = ~n20892 & ~n21510;
  assign n21512 = ~n20889 & ~n21511;
  assign n21513 = ~n20874 & ~n21512;
  assign n21514 = ~n20871 & ~n21513;
  assign n21515 = ~n20856 & ~n21514;
  assign n21516 = ~n20853 & ~n21515;
  assign n21517 = ~n20838 & ~n21516;
  assign n21518 = n20838 & n21516;
  assign n21519 = ~n21517 & ~n21518;
  assign n21520 = n20856 & n21514;
  assign n21521 = ~n21515 & ~n21520;
  assign n21522 = n11727 & ~n13438;
  assign n21523 = n11055 & ~n13627;
  assign n21524 = n11715 & n13941;
  assign n21525 = ~n21523 & ~n21524;
  assign n21526 = ~n21522 & n21525;
  assign n21527 = ~n11057 & n21526;
  assign n21528 = ~n14028 & n21526;
  assign n21529 = ~n21527 & ~n21528;
  assign n21530 =  a[2]  & ~n21529;
  assign n21531 = ~ a[2]  & n21529;
  assign n21532 = ~n21530 & ~n21531;
  assign n21533 = n21521 & ~n21532;
  assign n21534 = n20874 & n21512;
  assign n21535 = ~n21513 & ~n21534;
  assign n21536 = n11727 & n13941;
  assign n21537 = n11055 & n13633;
  assign n21538 = n11715 & ~n13627;
  assign n21539 = ~n21537 & ~n21538;
  assign n21540 = ~n21536 & n21539;
  assign n21541 = ~n11057 & n21540;
  assign n21542 = ~n14136 & n21540;
  assign n21543 = ~n21541 & ~n21542;
  assign n21544 =  a[2]  & ~n21543;
  assign n21545 = ~ a[2]  & n21543;
  assign n21546 = ~n21544 & ~n21545;
  assign n21547 = n21535 & ~n21546;
  assign n21548 = n20892 & n21510;
  assign n21549 = ~n21511 & ~n21548;
  assign n21550 = n11727 & ~n13627;
  assign n21551 = n11055 & n13630;
  assign n21552 = n11715 & n13633;
  assign n21553 = ~n21551 & ~n21552;
  assign n21554 = ~n21550 & n21553;
  assign n21555 = ~n11057 & n21554;
  assign n21556 = n13654 & n21554;
  assign n21557 = ~n21555 & ~n21556;
  assign n21558 =  a[2]  & ~n21557;
  assign n21559 = ~ a[2]  & n21557;
  assign n21560 = ~n21558 & ~n21559;
  assign n21561 = n21549 & ~n21560;
  assign n21562 = n20910 & n21508;
  assign n21563 = ~n21509 & ~n21562;
  assign n21564 = n11727 & n13633;
  assign n21565 = n11055 & n13597;
  assign n21566 = n11715 & n13630;
  assign n21567 = ~n21565 & ~n21566;
  assign n21568 = ~n21564 & n21567;
  assign n21569 = ~n11057 & n21568;
  assign n21570 = ~n13929 & n21568;
  assign n21571 = ~n21569 & ~n21570;
  assign n21572 =  a[2]  & ~n21571;
  assign n21573 = ~ a[2]  & n21571;
  assign n21574 = ~n21572 & ~n21573;
  assign n21575 = n21563 & ~n21574;
  assign n21576 = n20928 & n21506;
  assign n21577 = ~n21507 & ~n21576;
  assign n21578 = n11727 & n13630;
  assign n21579 = n11055 & n13515;
  assign n21580 = n11715 & n13597;
  assign n21581 = ~n21579 & ~n21580;
  assign n21582 = ~n21578 & n21581;
  assign n21583 = ~n11057 & n21582;
  assign n21584 = ~n13976 & n21582;
  assign n21585 = ~n21583 & ~n21584;
  assign n21586 =  a[2]  & ~n21585;
  assign n21587 = ~ a[2]  & n21585;
  assign n21588 = ~n21586 & ~n21587;
  assign n21589 = n21577 & ~n21588;
  assign n21590 = n20946 & n21504;
  assign n21591 = ~n21505 & ~n21590;
  assign n21592 = n11727 & n13597;
  assign n21593 = n11055 & n13521;
  assign n21594 = n11715 & n13515;
  assign n21595 = ~n21593 & ~n21594;
  assign n21596 = ~n21592 & n21595;
  assign n21597 = ~n11057 & n21596;
  assign n21598 = n13612 & n21596;
  assign n21599 = ~n21597 & ~n21598;
  assign n21600 =  a[2]  & ~n21599;
  assign n21601 = ~ a[2]  & n21599;
  assign n21602 = ~n21600 & ~n21601;
  assign n21603 = n21591 & ~n21602;
  assign n21604 = n20964 & n21502;
  assign n21605 = ~n21503 & ~n21604;
  assign n21606 = n11727 & n13515;
  assign n21607 = n11055 & n13518;
  assign n21608 = n11715 & n13521;
  assign n21609 = ~n21607 & ~n21608;
  assign n21610 = ~n21606 & n21609;
  assign n21611 = ~n11057 & n21610;
  assign n21612 = ~n13541 & n21610;
  assign n21613 = ~n21611 & ~n21612;
  assign n21614 =  a[2]  & ~n21613;
  assign n21615 = ~ a[2]  & n21613;
  assign n21616 = ~n21614 & ~n21615;
  assign n21617 = n21605 & ~n21616;
  assign n21618 = n20982 & n21500;
  assign n21619 = ~n21501 & ~n21618;
  assign n21620 = n11727 & n13521;
  assign n21621 = n11055 & n13491;
  assign n21622 = n11715 & n13518;
  assign n21623 = ~n21621 & ~n21622;
  assign n21624 = ~n21620 & n21623;
  assign n21625 = ~n11057 & n21624;
  assign n21626 = n13909 & n21624;
  assign n21627 = ~n21625 & ~n21626;
  assign n21628 =  a[2]  & ~n21627;
  assign n21629 = ~ a[2]  & n21627;
  assign n21630 = ~n21628 & ~n21629;
  assign n21631 = n21619 & ~n21630;
  assign n21632 = n21000 & n21498;
  assign n21633 = ~n21499 & ~n21632;
  assign n21634 = n11727 & n13518;
  assign n21635 = n11055 & n12889;
  assign n21636 = n11715 & n13491;
  assign n21637 = ~n21635 & ~n21636;
  assign n21638 = ~n21634 & n21637;
  assign n21639 = ~n11057 & n21638;
  assign n21640 = ~n13584 & n21638;
  assign n21641 = ~n21639 & ~n21640;
  assign n21642 =  a[2]  & ~n21641;
  assign n21643 = ~ a[2]  & n21641;
  assign n21644 = ~n21642 & ~n21643;
  assign n21645 = n21633 & ~n21644;
  assign n21646 = n21494 & ~n21496;
  assign n21647 = ~n21497 & ~n21646;
  assign n21648 = n21479 & ~n21481;
  assign n21649 = ~n21482 & ~n21648;
  assign n21650 = n21459 & ~n21461;
  assign n21651 = ~n21462 & ~n21650;
  assign n21652 = n21439 & ~n21441;
  assign n21653 = ~n21442 & ~n21652;
  assign n21654 = n21417 & ~n21419;
  assign n21655 = ~n21420 & ~n21654;
  assign n21656 = ~n21388 & n21399;
  assign n21657 = ~n21400 & ~n21656;
  assign n21658 = ~n11794 & ~n12581;
  assign n21659 = n11796 & ~n16094;
  assign n21660 = n11727 & n12574;
  assign n21661 = n11055 & ~n12581;
  assign n21662 = n11715 & n12577;
  assign n21663 = ~n21661 & ~n21662;
  assign n21664 = ~n21660 & n21663;
  assign n21665 =  a[2]  & ~n21664;
  assign n21666 = n11796 & ~n16085;
  assign n21667 = n11805 & ~n12581;
  assign n21668 = n11807 & n12577;
  assign n21669 =  a[2]  & ~n21668;
  assign n21670 = ~n21667 & n21669;
  assign n21671 = ~n21666 & n21670;
  assign n21672 = ~n21665 & n21671;
  assign n21673 = ~n21659 & n21672;
  assign n21674 = ~n21658 & n21673;
  assign n21675 = n21386 & n21674;
  assign n21676 = ~n21386 & ~n21674;
  assign n21677 = n11727 & n12571;
  assign n21678 = n11055 & n12577;
  assign n21679 = n11715 & n12574;
  assign n21680 = ~n21678 & ~n21679;
  assign n21681 = ~n21677 & n21680;
  assign n21682 = n11057 & n16013;
  assign n21683 = n21681 & ~n21682;
  assign n21684 = ~ a[2]  & ~n21683;
  assign n21685 =  a[2]  & n21683;
  assign n21686 = ~n21684 & ~n21685;
  assign n21687 = ~n21676 & ~n21686;
  assign n21688 = ~n21675 & ~n21687;
  assign n21689 = n11727 & n12567;
  assign n21690 = n11055 & n12574;
  assign n21691 = n11715 & n12571;
  assign n21692 = ~n21690 & ~n21691;
  assign n21693 = ~n21689 & n21692;
  assign n21694 = ~n11057 & n21693;
  assign n21695 = ~n15989 & n21693;
  assign n21696 = ~n21694 & ~n21695;
  assign n21697 =  a[2]  & ~n21696;
  assign n21698 = ~ a[2]  & n21696;
  assign n21699 = ~n21697 & ~n21698;
  assign n21700 = n21688 & n21699;
  assign n21701 = n21385 & ~n21387;
  assign n21702 = ~n21388 & ~n21701;
  assign n21703 = ~n21700 & n21702;
  assign n21704 = ~n21688 & ~n21699;
  assign n21705 = ~n21703 & ~n21704;
  assign n21706 = n21657 & ~n21705;
  assign n21707 = ~n21657 & n21705;
  assign n21708 = n11727 & n12564;
  assign n21709 = n11055 & n12571;
  assign n21710 = n11715 & n12567;
  assign n21711 = ~n21709 & ~n21710;
  assign n21712 = ~n21708 & n21711;
  assign n21713 = n11057 & ~n15944;
  assign n21714 = n21712 & ~n21713;
  assign n21715 = ~ a[2]  & ~n21714;
  assign n21716 =  a[2]  & n21714;
  assign n21717 = ~n21715 & ~n21716;
  assign n21718 = ~n21707 & ~n21717;
  assign n21719 = ~n21706 & ~n21718;
  assign n21720 = n11727 & n12561;
  assign n21721 = n11055 & n12567;
  assign n21722 = n11715 & n12564;
  assign n21723 = ~n21721 & ~n21722;
  assign n21724 = ~n21720 & n21723;
  assign n21725 = ~n11057 & n21724;
  assign n21726 = n15905 & n21724;
  assign n21727 = ~n21725 & ~n21726;
  assign n21728 =  a[2]  & ~n21727;
  assign n21729 = ~ a[2]  & n21727;
  assign n21730 = ~n21728 & ~n21729;
  assign n21731 = ~n21719 & ~n21730;
  assign n21732 = n21719 & n21730;
  assign n21733 = n21404 & n21415;
  assign n21734 = ~n21416 & ~n21733;
  assign n21735 = ~n21732 & n21734;
  assign n21736 = ~n21731 & ~n21735;
  assign n21737 = n21655 & ~n21736;
  assign n21738 = ~n21655 & n21736;
  assign n21739 = n11727 & n12558;
  assign n21740 = n11055 & n12564;
  assign n21741 = n11715 & n12561;
  assign n21742 = ~n21740 & ~n21741;
  assign n21743 = ~n21739 & n21742;
  assign n21744 = n11057 & n15847;
  assign n21745 = n21743 & ~n21744;
  assign n21746 = ~ a[2]  & ~n21745;
  assign n21747 =  a[2]  & n21745;
  assign n21748 = ~n21746 & ~n21747;
  assign n21749 = ~n21738 & ~n21748;
  assign n21750 = ~n21737 & ~n21749;
  assign n21751 = n11727 & n12555;
  assign n21752 = n11055 & n12561;
  assign n21753 = n11715 & n12558;
  assign n21754 = ~n21752 & ~n21753;
  assign n21755 = ~n21751 & n21754;
  assign n21756 = ~n11057 & n21755;
  assign n21757 = n15816 & n21755;
  assign n21758 = ~n21756 & ~n21757;
  assign n21759 =  a[2]  & ~n21758;
  assign n21760 = ~ a[2]  & n21758;
  assign n21761 = ~n21759 & ~n21760;
  assign n21762 = n21750 & n21761;
  assign n21763 = n21362 & n21421;
  assign n21764 = ~n21422 & ~n21763;
  assign n21765 = ~n21762 & n21764;
  assign n21766 = ~n21750 & ~n21761;
  assign n21767 = ~n21765 & ~n21766;
  assign n21768 = n11727 & n12552;
  assign n21769 = n11055 & n12558;
  assign n21770 = n11715 & n12555;
  assign n21771 = ~n21769 & ~n21770;
  assign n21772 = ~n21768 & n21771;
  assign n21773 = ~n11057 & n21772;
  assign n21774 = n15791 & n21772;
  assign n21775 = ~n21773 & ~n21774;
  assign n21776 =  a[2]  & ~n21775;
  assign n21777 = ~ a[2]  & n21775;
  assign n21778 = ~n21776 & ~n21777;
  assign n21779 = n21767 & n21778;
  assign n21780 = n21423 & ~n21425;
  assign n21781 = ~n21426 & ~n21780;
  assign n21782 = ~n21779 & n21781;
  assign n21783 = ~n21767 & ~n21778;
  assign n21784 = ~n21782 & ~n21783;
  assign n21785 = n11727 & n12549;
  assign n21786 = n11055 & n12555;
  assign n21787 = n11715 & n12552;
  assign n21788 = ~n21786 & ~n21787;
  assign n21789 = ~n21785 & n21788;
  assign n21790 = ~n11057 & n21789;
  assign n21791 = ~n15764 & n21789;
  assign n21792 = ~n21790 & ~n21791;
  assign n21793 =  a[2]  & ~n21792;
  assign n21794 = ~ a[2]  & n21792;
  assign n21795 = ~n21793 & ~n21794;
  assign n21796 = n21784 & n21795;
  assign n21797 = n21330 & n21427;
  assign n21798 = ~n21428 & ~n21797;
  assign n21799 = ~n21796 & n21798;
  assign n21800 = ~n21784 & ~n21795;
  assign n21801 = ~n21799 & ~n21800;
  assign n21802 = n21429 & ~n21431;
  assign n21803 = ~n21430 & n21802;
  assign n21804 = ~n21433 & ~n21803;
  assign n21805 = ~n21801 & n21804;
  assign n21806 = n21801 & ~n21804;
  assign n21807 = n11727 & n12546;
  assign n21808 = n11055 & n12552;
  assign n21809 = n11715 & n12549;
  assign n21810 = ~n21808 & ~n21809;
  assign n21811 = ~n21807 & n21810;
  assign n21812 = n11057 & ~n15356;
  assign n21813 = n21811 & ~n21812;
  assign n21814 = ~ a[2]  & ~n21813;
  assign n21815 =  a[2]  & n21813;
  assign n21816 = ~n21814 & ~n21815;
  assign n21817 = ~n21806 & ~n21816;
  assign n21818 = ~n21805 & ~n21817;
  assign n21819 = n21434 & ~n21436;
  assign n21820 = ~n21435 & n21819;
  assign n21821 = ~n21438 & ~n21820;
  assign n21822 = ~n21818 & n21821;
  assign n21823 = n21818 & ~n21821;
  assign n21824 = n11727 & n12543;
  assign n21825 = n11055 & n12549;
  assign n21826 = n11715 & n12546;
  assign n21827 = ~n21825 & ~n21826;
  assign n21828 = ~n21824 & n21827;
  assign n21829 = n11057 & n15724;
  assign n21830 = n21828 & ~n21829;
  assign n21831 = ~ a[2]  & ~n21830;
  assign n21832 =  a[2]  & n21830;
  assign n21833 = ~n21831 & ~n21832;
  assign n21834 = ~n21823 & ~n21833;
  assign n21835 = ~n21822 & ~n21834;
  assign n21836 = n21653 & ~n21835;
  assign n21837 = ~n21653 & n21835;
  assign n21838 = n11727 & n12540;
  assign n21839 = n11055 & n12546;
  assign n21840 = n11715 & n12543;
  assign n21841 = ~n21839 & ~n21840;
  assign n21842 = ~n21838 & n21841;
  assign n21843 = n11057 & ~n15708;
  assign n21844 = n21842 & ~n21843;
  assign n21845 = ~ a[2]  & ~n21844;
  assign n21846 =  a[2]  & n21844;
  assign n21847 = ~n21845 & ~n21846;
  assign n21848 = ~n21837 & ~n21847;
  assign n21849 = ~n21836 & ~n21848;
  assign n21850 = n11727 & n12537;
  assign n21851 = n11055 & n12543;
  assign n21852 = n11715 & n12540;
  assign n21853 = ~n21851 & ~n21852;
  assign n21854 = ~n21850 & n21853;
  assign n21855 = ~n11057 & n21854;
  assign n21856 = n15385 & n21854;
  assign n21857 = ~n21855 & ~n21856;
  assign n21858 =  a[2]  & ~n21857;
  assign n21859 = ~ a[2]  & n21857;
  assign n21860 = ~n21858 & ~n21859;
  assign n21861 = n21849 & n21860;
  assign n21862 = n21271 & n21443;
  assign n21863 = ~n21444 & ~n21862;
  assign n21864 = ~n21861 & n21863;
  assign n21865 = ~n21849 & ~n21860;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = n11727 & n12534;
  assign n21868 = n11055 & n12540;
  assign n21869 = n11715 & n12537;
  assign n21870 = ~n21868 & ~n21869;
  assign n21871 = ~n21867 & n21870;
  assign n21872 = ~n11057 & n21871;
  assign n21873 = n15096 & n21871;
  assign n21874 = ~n21872 & ~n21873;
  assign n21875 =  a[2]  & ~n21874;
  assign n21876 = ~ a[2]  & n21874;
  assign n21877 = ~n21875 & ~n21876;
  assign n21878 = n21866 & n21877;
  assign n21879 = n21253 & n21445;
  assign n21880 = ~n21446 & ~n21879;
  assign n21881 = ~n21878 & n21880;
  assign n21882 = ~n21866 & ~n21877;
  assign n21883 = ~n21881 & ~n21882;
  assign n21884 = n11727 & n12531;
  assign n21885 = n11055 & n12537;
  assign n21886 = n11715 & n12534;
  assign n21887 = ~n21885 & ~n21886;
  assign n21888 = ~n21884 & n21887;
  assign n21889 = ~n11057 & n21888;
  assign n21890 = ~n15255 & n21888;
  assign n21891 = ~n21889 & ~n21890;
  assign n21892 =  a[2]  & ~n21891;
  assign n21893 = ~ a[2]  & n21891;
  assign n21894 = ~n21892 & ~n21893;
  assign n21895 = n21883 & n21894;
  assign n21896 = n21235 & n21447;
  assign n21897 = ~n21448 & ~n21896;
  assign n21898 = ~n21895 & n21897;
  assign n21899 = ~n21883 & ~n21894;
  assign n21900 = ~n21898 & ~n21899;
  assign n21901 = n21449 & ~n21451;
  assign n21902 = ~n21450 & n21901;
  assign n21903 = ~n21453 & ~n21902;
  assign n21904 = ~n21900 & n21903;
  assign n21905 = n21900 & ~n21903;
  assign n21906 = n11727 & n12528;
  assign n21907 = n11055 & n12534;
  assign n21908 = n11715 & n12531;
  assign n21909 = ~n21907 & ~n21908;
  assign n21910 = ~n21906 & n21909;
  assign n21911 = n11057 & ~n15003;
  assign n21912 = n21910 & ~n21911;
  assign n21913 = ~ a[2]  & ~n21912;
  assign n21914 =  a[2]  & n21912;
  assign n21915 = ~n21913 & ~n21914;
  assign n21916 = ~n21905 & ~n21915;
  assign n21917 = ~n21904 & ~n21916;
  assign n21918 = n21454 & ~n21456;
  assign n21919 = ~n21455 & n21918;
  assign n21920 = ~n21458 & ~n21919;
  assign n21921 = ~n21917 & n21920;
  assign n21922 = n21917 & ~n21920;
  assign n21923 = n11727 & n12525;
  assign n21924 = n11055 & n12531;
  assign n21925 = n11715 & n12528;
  assign n21926 = ~n21924 & ~n21925;
  assign n21927 = ~n21923 & n21926;
  assign n21928 = n11057 & n14608;
  assign n21929 = n21927 & ~n21928;
  assign n21930 = ~ a[2]  & ~n21929;
  assign n21931 =  a[2]  & n21929;
  assign n21932 = ~n21930 & ~n21931;
  assign n21933 = ~n21922 & ~n21932;
  assign n21934 = ~n21921 & ~n21933;
  assign n21935 = n21651 & ~n21934;
  assign n21936 = ~n21651 & n21934;
  assign n21937 = n11727 & n12522;
  assign n21938 = n11055 & n12528;
  assign n21939 = n11715 & n12525;
  assign n21940 = ~n21938 & ~n21939;
  assign n21941 = ~n21937 & n21940;
  assign n21942 = n11057 & n14837;
  assign n21943 = n21941 & ~n21942;
  assign n21944 = ~ a[2]  & ~n21943;
  assign n21945 =  a[2]  & n21943;
  assign n21946 = ~n21944 & ~n21945;
  assign n21947 = ~n21936 & ~n21946;
  assign n21948 = ~n21935 & ~n21947;
  assign n21949 = n11727 & n12519;
  assign n21950 = n11055 & n12525;
  assign n21951 = n11715 & n12522;
  assign n21952 = ~n21950 & ~n21951;
  assign n21953 = ~n21949 & n21952;
  assign n21954 = ~n11057 & n21953;
  assign n21955 = ~n14454 & n21953;
  assign n21956 = ~n21954 & ~n21955;
  assign n21957 =  a[2]  & ~n21956;
  assign n21958 = ~ a[2]  & n21956;
  assign n21959 = ~n21957 & ~n21958;
  assign n21960 = n21948 & n21959;
  assign n21961 = n21176 & n21463;
  assign n21962 = ~n21464 & ~n21961;
  assign n21963 = ~n21960 & n21962;
  assign n21964 = ~n21948 & ~n21959;
  assign n21965 = ~n21963 & ~n21964;
  assign n21966 = n11727 & n12516;
  assign n21967 = n11055 & n12522;
  assign n21968 = n11715 & n12519;
  assign n21969 = ~n21967 & ~n21968;
  assign n21970 = ~n21966 & n21969;
  assign n21971 = ~n11057 & n21970;
  assign n21972 = n14443 & n21970;
  assign n21973 = ~n21971 & ~n21972;
  assign n21974 =  a[2]  & ~n21973;
  assign n21975 = ~ a[2]  & n21973;
  assign n21976 = ~n21974 & ~n21975;
  assign n21977 = n21965 & n21976;
  assign n21978 = n21158 & n21465;
  assign n21979 = ~n21466 & ~n21978;
  assign n21980 = ~n21977 & n21979;
  assign n21981 = ~n21965 & ~n21976;
  assign n21982 = ~n21980 & ~n21981;
  assign n21983 = n11727 & n12511;
  assign n21984 = n11055 & n12519;
  assign n21985 = n11715 & n12516;
  assign n21986 = ~n21984 & ~n21985;
  assign n21987 = ~n21983 & n21986;
  assign n21988 = ~n11057 & n21987;
  assign n21989 = n14233 & n21987;
  assign n21990 = ~n21988 & ~n21989;
  assign n21991 =  a[2]  & ~n21990;
  assign n21992 = ~ a[2]  & n21990;
  assign n21993 = ~n21991 & ~n21992;
  assign n21994 = n21982 & n21993;
  assign n21995 = n21140 & n21467;
  assign n21996 = ~n21468 & ~n21995;
  assign n21997 = ~n21994 & n21996;
  assign n21998 = ~n21982 & ~n21993;
  assign n21999 = ~n21997 & ~n21998;
  assign n22000 = n21469 & ~n21471;
  assign n22001 = ~n21470 & n22000;
  assign n22002 = ~n21473 & ~n22001;
  assign n22003 = ~n21999 & n22002;
  assign n22004 = n21999 & ~n22002;
  assign n22005 = n11727 & n12513;
  assign n22006 = n11055 & n12516;
  assign n22007 = n11715 & n12511;
  assign n22008 = ~n22006 & ~n22007;
  assign n22009 = ~n22005 & n22008;
  assign n22010 = n11057 & n14177;
  assign n22011 = n22009 & ~n22010;
  assign n22012 = ~ a[2]  & ~n22011;
  assign n22013 =  a[2]  & n22011;
  assign n22014 = ~n22012 & ~n22013;
  assign n22015 = ~n22004 & ~n22014;
  assign n22016 = ~n22003 & ~n22015;
  assign n22017 = n21474 & ~n21476;
  assign n22018 = ~n21475 & n22017;
  assign n22019 = ~n21478 & ~n22018;
  assign n22020 = ~n22016 & n22019;
  assign n22021 = n22016 & ~n22019;
  assign n22022 = n11727 & n12508;
  assign n22023 = n11055 & n12511;
  assign n22024 = n11715 & n12513;
  assign n22025 = ~n22023 & ~n22024;
  assign n22026 = ~n22022 & n22025;
  assign n22027 = n11057 & n13863;
  assign n22028 = n22026 & ~n22027;
  assign n22029 = ~ a[2]  & ~n22028;
  assign n22030 =  a[2]  & n22028;
  assign n22031 = ~n22029 & ~n22030;
  assign n22032 = ~n22021 & ~n22031;
  assign n22033 = ~n22020 & ~n22032;
  assign n22034 = n21649 & ~n22033;
  assign n22035 = ~n21649 & n22033;
  assign n22036 = n11727 & n12505;
  assign n22037 = n11055 & n12513;
  assign n22038 = n11715 & n12508;
  assign n22039 = ~n22037 & ~n22038;
  assign n22040 = ~n22036 & n22039;
  assign n22041 = n11057 & ~n14051;
  assign n22042 = n22040 & ~n22041;
  assign n22043 = ~ a[2]  & ~n22042;
  assign n22044 =  a[2]  & n22042;
  assign n22045 = ~n22043 & ~n22044;
  assign n22046 = ~n22035 & ~n22045;
  assign n22047 = ~n22034 & ~n22046;
  assign n22048 = n11727 & n12370;
  assign n22049 = n11055 & n12508;
  assign n22050 = n11715 & n12505;
  assign n22051 = ~n22049 & ~n22050;
  assign n22052 = ~n22048 & n22051;
  assign n22053 = ~n11057 & n22052;
  assign n22054 = n13748 & n22052;
  assign n22055 = ~n22053 & ~n22054;
  assign n22056 =  a[2]  & ~n22055;
  assign n22057 = ~ a[2]  & n22055;
  assign n22058 = ~n22056 & ~n22057;
  assign n22059 = n22047 & n22058;
  assign n22060 = n21081 & n21483;
  assign n22061 = ~n21484 & ~n22060;
  assign n22062 = ~n22059 & n22061;
  assign n22063 = ~n22047 & ~n22058;
  assign n22064 = ~n22062 & ~n22063;
  assign n22065 = n11727 & n12502;
  assign n22066 = n11055 & n12505;
  assign n22067 = n11715 & n12370;
  assign n22068 = ~n22066 & ~n22067;
  assign n22069 = ~n22065 & n22068;
  assign n22070 = ~n11057 & n22069;
  assign n22071 = n13736 & n22069;
  assign n22072 = ~n22070 & ~n22071;
  assign n22073 =  a[2]  & ~n22072;
  assign n22074 = ~ a[2]  & n22072;
  assign n22075 = ~n22073 & ~n22074;
  assign n22076 = n22064 & n22075;
  assign n22077 = n21063 & n21485;
  assign n22078 = ~n21486 & ~n22077;
  assign n22079 = ~n22076 & n22078;
  assign n22080 = ~n22064 & ~n22075;
  assign n22081 = ~n22079 & ~n22080;
  assign n22082 = n11727 & n12769;
  assign n22083 = n11055 & n12370;
  assign n22084 = n11715 & n12502;
  assign n22085 = ~n22083 & ~n22084;
  assign n22086 = ~n22082 & n22085;
  assign n22087 = ~n11057 & n22086;
  assign n22088 = ~n12999 & n22086;
  assign n22089 = ~n22087 & ~n22088;
  assign n22090 =  a[2]  & ~n22089;
  assign n22091 = ~ a[2]  & n22089;
  assign n22092 = ~n22090 & ~n22091;
  assign n22093 = n22081 & n22092;
  assign n22094 = n21045 & n21487;
  assign n22095 = ~n21488 & ~n22094;
  assign n22096 = ~n22093 & n22095;
  assign n22097 = ~n22081 & ~n22092;
  assign n22098 = ~n22096 & ~n22097;
  assign n22099 = n21489 & ~n21491;
  assign n22100 = ~n21490 & n22099;
  assign n22101 = ~n21493 & ~n22100;
  assign n22102 = ~n22098 & n22101;
  assign n22103 = n22098 & ~n22101;
  assign n22104 = n11727 & n12889;
  assign n22105 = n11055 & n12502;
  assign n22106 = n11715 & n12769;
  assign n22107 = ~n22105 & ~n22106;
  assign n22108 = ~n22104 & n22107;
  assign n22109 = n11057 & n12895;
  assign n22110 = n22108 & ~n22109;
  assign n22111 = ~ a[2]  & ~n22110;
  assign n22112 =  a[2]  & n22110;
  assign n22113 = ~n22111 & ~n22112;
  assign n22114 = ~n22103 & ~n22113;
  assign n22115 = ~n22102 & ~n22114;
  assign n22116 = n21647 & ~n22115;
  assign n22117 = ~n21647 & n22115;
  assign n22118 = n11727 & n13491;
  assign n22119 = n11055 & n12769;
  assign n22120 = n11715 & n12889;
  assign n22121 = ~n22119 & ~n22120;
  assign n22122 = ~n22118 & n22121;
  assign n22123 = n11057 & ~n13503;
  assign n22124 = n22122 & ~n22123;
  assign n22125 = ~ a[2]  & ~n22124;
  assign n22126 =  a[2]  & n22124;
  assign n22127 = ~n22125 & ~n22126;
  assign n22128 = ~n22117 & ~n22127;
  assign n22129 = ~n22116 & ~n22128;
  assign n22130 = n21633 & ~n21645;
  assign n22131 = ~n21644 & ~n21645;
  assign n22132 = ~n22130 & ~n22131;
  assign n22133 = ~n22129 & ~n22132;
  assign n22134 = ~n21645 & ~n22133;
  assign n22135 = ~n21619 & n21630;
  assign n22136 = ~n21631 & ~n22135;
  assign n22137 = ~n22134 & n22136;
  assign n22138 = ~n21631 & ~n22137;
  assign n22139 = ~n21605 & n21616;
  assign n22140 = ~n21617 & ~n22139;
  assign n22141 = ~n22138 & n22140;
  assign n22142 = ~n21617 & ~n22141;
  assign n22143 = ~n21591 & n21602;
  assign n22144 = ~n21603 & ~n22143;
  assign n22145 = ~n22142 & n22144;
  assign n22146 = ~n21603 & ~n22145;
  assign n22147 = ~n21577 & n21588;
  assign n22148 = ~n21589 & ~n22147;
  assign n22149 = ~n22146 & n22148;
  assign n22150 = ~n21589 & ~n22149;
  assign n22151 = ~n21563 & n21574;
  assign n22152 = ~n21575 & ~n22151;
  assign n22153 = ~n22150 & n22152;
  assign n22154 = ~n21575 & ~n22153;
  assign n22155 = ~n21549 & n21560;
  assign n22156 = ~n21561 & ~n22155;
  assign n22157 = ~n22154 & n22156;
  assign n22158 = ~n21561 & ~n22157;
  assign n22159 = ~n21535 & n21546;
  assign n22160 = ~n21547 & ~n22159;
  assign n22161 = ~n22158 & n22160;
  assign n22162 = ~n21547 & ~n22161;
  assign n22163 = ~n21521 & n21532;
  assign n22164 = ~n21533 & ~n22163;
  assign n22165 = ~n22162 & n22164;
  assign n22166 = ~n21533 & ~n22165;
  assign n22167 = n21519 & ~n22166;
  assign n22168 = ~n21517 & ~n22167;
  assign n22169 = n20835 & ~n22168;
  assign n22170 = ~n20833 & ~n22169;
  assign n22171 = n20800 & ~n22170;
  assign n22172 = ~n20798 & ~n22171;
  assign n22173 = n20145 & ~n22172;
  assign n22174 = ~n20143 & ~n22173;
  assign n22175 = n19516 & ~n19518;
  assign n22176 = ~n19519 & ~n22175;
  assign n22177 = ~n22174 & n22176;
  assign n22178 = ~n19519 & ~n22177;
  assign n22179 = ~n18946 & ~n22178;
  assign n22180 = ~n18943 & ~n22179;
  assign n22181 = n18396 & ~n22180;
  assign n22182 = ~n18394 & ~n22181;
  assign n22183 = n17892 & ~n17894;
  assign n22184 = ~n17895 & ~n22183;
  assign n22185 = ~n22182 & n22184;
  assign n22186 = ~n17895 & ~n22185;
  assign n22187 = ~n17428 & ~n22186;
  assign n22188 = ~n17425 & ~n22187;
  assign n22189 = n17001 & ~n22188;
  assign n22190 = ~n16999 & ~n22189;
  assign n22191 = n16604 & ~n16606;
  assign n22192 = ~n16607 & ~n22191;
  assign n22193 = ~n22190 & n22192;
  assign n22194 = ~n16607 & ~n22193;
  assign n22195 = ~n16443 & ~n22194;
  assign n22196 = ~n16440 & ~n22195;
  assign n22197 = n16272 & ~n22196;
  assign n22198 = ~n16270 & ~n22197;
  assign n22199 = n15650 & ~n15652;
  assign n22200 = ~n15653 & ~n22199;
  assign n22201 = ~n22198 & n22200;
  assign n22202 = ~n15653 & ~n22201;
  assign n22203 = ~n15508 & ~n22202;
  assign n22204 = ~n15505 & ~n22203;
  assign n22205 = n15203 & ~n22204;
  assign n22206 = ~n15201 & ~n22205;
  assign n22207 = n14950 & ~n14952;
  assign n22208 = ~n14953 & ~n22207;
  assign n22209 = ~n22206 & n22208;
  assign n22210 = ~n14953 & ~n22209;
  assign n22211 = ~n14809 & ~n22210;
  assign n22212 = ~n14806 & ~n22211;
  assign n22213 = n14696 & ~n22212;
  assign n22214 = ~n14694 & ~n22213;
  assign n22215 = n14321 & ~n14323;
  assign n22216 = ~n14324 & ~n22215;
  assign n22217 = ~n22214 & n22216;
  assign n22218 = ~n14324 & ~n22217;
  assign n22219 = ~n14154 & ~n22218;
  assign n22220 = ~n14151 & ~n22219;
  assign n22221 = n14039 & ~n22220;
  assign n22222 = ~n14037 & ~n22221;
  assign n22223 = ~n13957 & ~n13960;
  assign n22224 = ~n13621 & ~n13661;
  assign n22225 = n3884 & n13941;
  assign n22226 = n3967 & n13633;
  assign n22227 = n4046 & ~n13627;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = ~n22225 & n22228;
  assign n22230 = n4050 & n14136;
  assign n22231 = n22229 & ~n22230;
  assign n22232 =  a[26]  & ~n22231;
  assign n22233 =  a[26]  & ~n22232;
  assign n22234 = ~n22231 & ~n22232;
  assign n22235 = ~n22233 & ~n22234;
  assign n22236 = ~n22224 & ~n22235;
  assign n22237 = ~n22224 & ~n22236;
  assign n22238 = ~n22235 & ~n22236;
  assign n22239 = ~n22237 & ~n22238;
  assign n22240 = n75 & ~n13909;
  assign n22241 = n3020 & n13521;
  assign n22242 = n3023 & n13491;
  assign n22243 = n3028 & n13518;
  assign n22244 = ~n22242 & ~n22243;
  assign n22245 = ~n22241 & n22244;
  assign n22246 = ~n22240 & n22245;
  assign n22247 = ~n4533 & n13938;
  assign n22248 = ~n4536 & n22247;
  assign n22249 = ~n13438 & ~n22248;
  assign n22250 =  a[23]  & ~n22249;
  assign n22251 = ~ a[23]  & n22249;
  assign n22252 = ~n22250 & ~n22251;
  assign n22253 = n303 & n3042;
  assign n22254 = n6567 & n22253;
  assign n22255 = n4827 & n22254;
  assign n22256 = n16031 & n22255;
  assign n22257 = n13787 & n22256;
  assign n22258 = n14534 & n22257;
  assign n22259 = n774 & n22258;
  assign n22260 = n471 & n22259;
  assign n22261 = n3733 & n22260;
  assign n22262 = n1269 & n22261;
  assign n22263 = ~n847 & n22262;
  assign n22264 = ~n367 & n22263;
  assign n22265 = ~n226 & n22264;
  assign n22266 = ~n306 & n22265;
  assign n22267 = ~n158 & n22266;
  assign n22268 = ~n270 & n22267;
  assign n22269 = n13574 & n22268;
  assign n22270 = ~n13574 & ~n22268;
  assign n22271 = ~n22269 & ~n22270;
  assign n22272 = n22252 & n22271;
  assign n22273 = ~n22252 & ~n22271;
  assign n22274 = ~n22272 & ~n22273;
  assign n22275 = ~n13580 & n22274;
  assign n22276 = n13580 & ~n22274;
  assign n22277 = ~n22275 & ~n22276;
  assign n22278 = ~n22246 & n22277;
  assign n22279 = n22277 & ~n22278;
  assign n22280 = ~n22246 & ~n22278;
  assign n22281 = ~n22279 & ~n22280;
  assign n22282 = ~n13592 & ~n13618;
  assign n22283 = n22281 & n22282;
  assign n22284 = ~n22281 & ~n22282;
  assign n22285 = ~n22283 & ~n22284;
  assign n22286 = n3457 & n13630;
  assign n22287 = n3542 & n13515;
  assign n22288 = n3606 & n13597;
  assign n22289 = ~n22287 & ~n22288;
  assign n22290 = ~n22286 & n22289;
  assign n22291 = n3368 & n13976;
  assign n22292 = n22290 & ~n22291;
  assign n22293 =  a[29]  & ~n22292;
  assign n22294 =  a[29]  & ~n22293;
  assign n22295 = ~n22292 & ~n22293;
  assign n22296 = ~n22294 & ~n22295;
  assign n22297 = n22285 & ~n22296;
  assign n22298 = n22285 & ~n22297;
  assign n22299 = ~n22296 & ~n22297;
  assign n22300 = ~n22298 & ~n22299;
  assign n22301 = ~n22239 & n22300;
  assign n22302 = n22239 & ~n22300;
  assign n22303 = ~n22301 & ~n22302;
  assign n22304 = ~n22223 & ~n22303;
  assign n22305 = n22223 & n22303;
  assign n22306 = ~n22304 & ~n22305;
  assign n22307 = ~n22222 & n22306;
  assign n22308 = n22222 & ~n22306;
  assign n22309 = ~n22307 & ~n22308;
  assign n22310 = n71 & n22309;
  assign n22311 = n14154 & n22218;
  assign n22312 = ~n22219 & ~n22311;
  assign n22313 = n9867 & n22312;
  assign n22314 = ~n14039 & n22220;
  assign n22315 = ~n22221 & ~n22314;
  assign n22316 = n10434 & n22315;
  assign n22317 = ~n22313 & ~n22316;
  assign n22318 = ~n22310 & n22317;
  assign n22319 = n22214 & ~n22216;
  assign n22320 = ~n22217 & ~n22319;
  assign n22321 = n22312 & n22320;
  assign n22322 = ~n14696 & n22212;
  assign n22323 = ~n22213 & ~n22322;
  assign n22324 = n22320 & n22323;
  assign n22325 = n14809 & n22210;
  assign n22326 = ~n22211 & ~n22325;
  assign n22327 = n22323 & n22326;
  assign n22328 = n22206 & ~n22208;
  assign n22329 = ~n22209 & ~n22328;
  assign n22330 = n22326 & n22329;
  assign n22331 = ~n15203 & n22204;
  assign n22332 = ~n22205 & ~n22331;
  assign n22333 = n22329 & n22332;
  assign n22334 = n15508 & n22202;
  assign n22335 = ~n22203 & ~n22334;
  assign n22336 = n22332 & n22335;
  assign n22337 = n22198 & ~n22200;
  assign n22338 = ~n22201 & ~n22337;
  assign n22339 = n22335 & n22338;
  assign n22340 = ~n16272 & n22196;
  assign n22341 = ~n22197 & ~n22340;
  assign n22342 = n22338 & n22341;
  assign n22343 = n16443 & n22194;
  assign n22344 = ~n22195 & ~n22343;
  assign n22345 = n22341 & n22344;
  assign n22346 = n22190 & ~n22192;
  assign n22347 = ~n22193 & ~n22346;
  assign n22348 = n22344 & n22347;
  assign n22349 = ~n17001 & n22188;
  assign n22350 = ~n22189 & ~n22349;
  assign n22351 = n22347 & n22350;
  assign n22352 = n17428 & n22186;
  assign n22353 = ~n22187 & ~n22352;
  assign n22354 = n22350 & n22353;
  assign n22355 = n22182 & ~n22184;
  assign n22356 = ~n22185 & ~n22355;
  assign n22357 = n22353 & n22356;
  assign n22358 = ~n18396 & n22180;
  assign n22359 = ~n22181 & ~n22358;
  assign n22360 = n22356 & n22359;
  assign n22361 = n18946 & n22178;
  assign n22362 = ~n22179 & ~n22361;
  assign n22363 = n22359 & n22362;
  assign n22364 = n22174 & ~n22176;
  assign n22365 = ~n22177 & ~n22364;
  assign n22366 = n22362 & n22365;
  assign n22367 = ~n20145 & n22172;
  assign n22368 = ~n22173 & ~n22367;
  assign n22369 = n22365 & n22368;
  assign n22370 = ~n20800 & n22170;
  assign n22371 = ~n22171 & ~n22370;
  assign n22372 = n22368 & n22371;
  assign n22373 = ~n20835 & n22168;
  assign n22374 = ~n22169 & ~n22373;
  assign n22375 = n22371 & n22374;
  assign n22376 = ~n21519 & n22166;
  assign n22377 = ~n22167 & ~n22376;
  assign n22378 = n22374 & n22377;
  assign n22379 = n22162 & ~n22164;
  assign n22380 = ~n22165 & ~n22379;
  assign n22381 = n22377 & n22380;
  assign n22382 = ~n22377 & ~n22380;
  assign n22383 = n22158 & ~n22160;
  assign n22384 = ~n22161 & ~n22383;
  assign n22385 = n22380 & n22384;
  assign n22386 = n22154 & ~n22156;
  assign n22387 = ~n22157 & ~n22386;
  assign n22388 = n22384 & n22387;
  assign n22389 = n22150 & ~n22152;
  assign n22390 = ~n22153 & ~n22389;
  assign n22391 = n22387 & n22390;
  assign n22392 = n22146 & ~n22148;
  assign n22393 = ~n22149 & ~n22392;
  assign n22394 = n22390 & n22393;
  assign n22395 = n22142 & ~n22144;
  assign n22396 = ~n22145 & ~n22395;
  assign n22397 = n22393 & n22396;
  assign n22398 = n22138 & ~n22140;
  assign n22399 = ~n22141 & ~n22398;
  assign n22400 = n22396 & n22399;
  assign n22401 = n22134 & ~n22136;
  assign n22402 = ~n22137 & ~n22401;
  assign n22403 = n22399 & n22402;
  assign n22404 = ~n22129 & ~n22133;
  assign n22405 = ~n22132 & ~n22133;
  assign n22406 = ~n22404 & ~n22405;
  assign n22407 = n22402 & ~n22406;
  assign n22408 = ~n22399 & n22407;
  assign n22409 = ~n22403 & ~n22408;
  assign n22410 = ~n22396 & ~n22399;
  assign n22411 = ~n22400 & ~n22410;
  assign n22412 = ~n22409 & n22411;
  assign n22413 = ~n22400 & ~n22412;
  assign n22414 = ~n22393 & ~n22396;
  assign n22415 = ~n22397 & ~n22414;
  assign n22416 = ~n22413 & n22415;
  assign n22417 = ~n22397 & ~n22416;
  assign n22418 = ~n22390 & ~n22393;
  assign n22419 = ~n22394 & ~n22418;
  assign n22420 = ~n22417 & n22419;
  assign n22421 = ~n22394 & ~n22420;
  assign n22422 = ~n22387 & ~n22390;
  assign n22423 = ~n22391 & ~n22422;
  assign n22424 = ~n22421 & n22423;
  assign n22425 = ~n22391 & ~n22424;
  assign n22426 = ~n22384 & ~n22387;
  assign n22427 = ~n22388 & ~n22426;
  assign n22428 = ~n22425 & n22427;
  assign n22429 = ~n22388 & ~n22428;
  assign n22430 = ~n22380 & ~n22384;
  assign n22431 = ~n22385 & ~n22430;
  assign n22432 = ~n22429 & n22431;
  assign n22433 = ~n22385 & ~n22432;
  assign n22434 = ~n22381 & ~n22433;
  assign n22435 = ~n22382 & n22434;
  assign n22436 = ~n22381 & ~n22435;
  assign n22437 = ~n22374 & ~n22377;
  assign n22438 = ~n22378 & ~n22437;
  assign n22439 = ~n22436 & n22438;
  assign n22440 = ~n22378 & ~n22439;
  assign n22441 = ~n22371 & ~n22374;
  assign n22442 = ~n22375 & ~n22441;
  assign n22443 = ~n22440 & n22442;
  assign n22444 = ~n22375 & ~n22443;
  assign n22445 = ~n22368 & ~n22371;
  assign n22446 = ~n22372 & ~n22445;
  assign n22447 = ~n22444 & n22446;
  assign n22448 = ~n22372 & ~n22447;
  assign n22449 = ~n22365 & ~n22368;
  assign n22450 = ~n22448 & ~n22449;
  assign n22451 = ~n22369 & n22450;
  assign n22452 = ~n22369 & ~n22451;
  assign n22453 = ~n22362 & ~n22365;
  assign n22454 = ~n22452 & ~n22453;
  assign n22455 = ~n22366 & n22454;
  assign n22456 = ~n22366 & ~n22455;
  assign n22457 = ~n22359 & ~n22362;
  assign n22458 = ~n22363 & ~n22457;
  assign n22459 = ~n22456 & n22458;
  assign n22460 = ~n22363 & ~n22459;
  assign n22461 = ~n22356 & ~n22359;
  assign n22462 = ~n22460 & ~n22461;
  assign n22463 = ~n22360 & n22462;
  assign n22464 = ~n22360 & ~n22463;
  assign n22465 = ~n22353 & ~n22356;
  assign n22466 = ~n22464 & ~n22465;
  assign n22467 = ~n22357 & n22466;
  assign n22468 = ~n22357 & ~n22467;
  assign n22469 = ~n22350 & ~n22353;
  assign n22470 = ~n22354 & ~n22469;
  assign n22471 = ~n22468 & n22470;
  assign n22472 = ~n22354 & ~n22471;
  assign n22473 = ~n22347 & ~n22350;
  assign n22474 = ~n22472 & ~n22473;
  assign n22475 = ~n22351 & n22474;
  assign n22476 = ~n22351 & ~n22475;
  assign n22477 = ~n22344 & ~n22347;
  assign n22478 = ~n22476 & ~n22477;
  assign n22479 = ~n22348 & n22478;
  assign n22480 = ~n22348 & ~n22479;
  assign n22481 = ~n22341 & ~n22344;
  assign n22482 = ~n22345 & ~n22481;
  assign n22483 = ~n22480 & n22482;
  assign n22484 = ~n22345 & ~n22483;
  assign n22485 = ~n22338 & ~n22341;
  assign n22486 = ~n22484 & ~n22485;
  assign n22487 = ~n22342 & n22486;
  assign n22488 = ~n22342 & ~n22487;
  assign n22489 = ~n22335 & ~n22338;
  assign n22490 = ~n22488 & ~n22489;
  assign n22491 = ~n22339 & n22490;
  assign n22492 = ~n22339 & ~n22491;
  assign n22493 = ~n22332 & ~n22335;
  assign n22494 = ~n22336 & ~n22493;
  assign n22495 = ~n22492 & n22494;
  assign n22496 = ~n22336 & ~n22495;
  assign n22497 = ~n22329 & ~n22332;
  assign n22498 = ~n22496 & ~n22497;
  assign n22499 = ~n22333 & n22498;
  assign n22500 = ~n22333 & ~n22499;
  assign n22501 = ~n22326 & ~n22329;
  assign n22502 = ~n22500 & ~n22501;
  assign n22503 = ~n22330 & n22502;
  assign n22504 = ~n22330 & ~n22503;
  assign n22505 = ~n22323 & ~n22326;
  assign n22506 = ~n22327 & ~n22505;
  assign n22507 = ~n22504 & n22506;
  assign n22508 = ~n22327 & ~n22507;
  assign n22509 = ~n22320 & ~n22323;
  assign n22510 = ~n22508 & ~n22509;
  assign n22511 = ~n22324 & n22510;
  assign n22512 = ~n22324 & ~n22511;
  assign n22513 = ~n22312 & ~n22320;
  assign n22514 = ~n22512 & ~n22513;
  assign n22515 = ~n22321 & n22514;
  assign n22516 = ~n22321 & ~n22515;
  assign n22517 = ~n22312 & ~n22315;
  assign n22518 = n22312 & n22315;
  assign n22519 = ~n22517 & ~n22518;
  assign n22520 = ~n22516 & n22519;
  assign n22521 = ~n22518 & ~n22520;
  assign n22522 = n22309 & n22315;
  assign n22523 = ~n22309 & ~n22315;
  assign n22524 = ~n22521 & ~n22523;
  assign n22525 = ~n22522 & n22524;
  assign n22526 = ~n22521 & ~n22525;
  assign n22527 = ~n22522 & ~n22525;
  assign n22528 = ~n22523 & n22527;
  assign n22529 = ~n22526 & ~n22528;
  assign n22530 = n9870 & ~n22529;
  assign n22531 = n22318 & ~n22530;
  assign n22532 =  a[5]  & ~n22531;
  assign n22533 = ~n22531 & ~n22532;
  assign n22534 =  a[5]  & ~n22532;
  assign n22535 = ~n22533 & ~n22534;
  assign n22536 = n7983 & n22332;
  assign n22537 = n7291 & n22338;
  assign n22538 = n7632 & n22335;
  assign n22539 = ~n22537 & ~n22538;
  assign n22540 = ~n22536 & n22539;
  assign n22541 = n22492 & ~n22494;
  assign n22542 = ~n22495 & ~n22541;
  assign n22543 = n7294 & n22542;
  assign n22544 = n22540 & ~n22543;
  assign n22545 =  a[11]  & ~n22544;
  assign n22546 = ~n22544 & ~n22545;
  assign n22547 =  a[11]  & ~n22545;
  assign n22548 = ~n22546 & ~n22547;
  assign n22549 = n6233 & n22353;
  assign n22550 = n5663 & n22359;
  assign n22551 = n5939 & n22356;
  assign n22552 = ~n22550 & ~n22551;
  assign n22553 = ~n22549 & n22552;
  assign n22554 = ~n22464 & ~n22467;
  assign n22555 = ~n22465 & n22468;
  assign n22556 = ~n22554 & ~n22555;
  assign n22557 = n5666 & ~n22556;
  assign n22558 = n22553 & ~n22557;
  assign n22559 =  a[17]  & ~n22558;
  assign n22560 = ~n22558 & ~n22559;
  assign n22561 =  a[17]  & ~n22559;
  assign n22562 = ~n22560 & ~n22561;
  assign n22563 = n4694 & n22374;
  assign n22564 = n4533 & n22380;
  assign n22565 = n4604 & n22377;
  assign n22566 = ~n22564 & ~n22565;
  assign n22567 = ~n22563 & n22566;
  assign n22568 = n22436 & ~n22438;
  assign n22569 = ~n22439 & ~n22568;
  assign n22570 = n4536 & n22569;
  assign n22571 = n22567 & ~n22570;
  assign n22572 =  a[23]  & ~n22571;
  assign n22573 = ~n22571 & ~n22572;
  assign n22574 =  a[23]  & ~n22572;
  assign n22575 = ~n22573 & ~n22574;
  assign n22576 = n3884 & n22387;
  assign n22577 = n3967 & n22393;
  assign n22578 = n4046 & n22390;
  assign n22579 = ~n22577 & ~n22578;
  assign n22580 = ~n22576 & n22579;
  assign n22581 = n22421 & ~n22423;
  assign n22582 = ~n22424 & ~n22581;
  assign n22583 = n4050 & n22582;
  assign n22584 = n22580 & ~n22583;
  assign n22585 =  a[26]  & ~n22584;
  assign n22586 = ~n22584 & ~n22585;
  assign n22587 =  a[26]  & ~n22585;
  assign n22588 = ~n22586 & ~n22587;
  assign n22589 = n3457 & n22396;
  assign n22590 = n3542 & n22402;
  assign n22591 = n3606 & n22399;
  assign n22592 = ~n22590 & ~n22591;
  assign n22593 = ~n22589 & n22592;
  assign n22594 = n22409 & ~n22411;
  assign n22595 = ~n22412 & ~n22594;
  assign n22596 = n3368 & n22595;
  assign n22597 = n22593 & ~n22596;
  assign n22598 =  a[29]  & ~n22597;
  assign n22599 = ~n22597 & ~n22598;
  assign n22600 =  a[29]  & ~n22598;
  assign n22601 = ~n22599 & ~n22600;
  assign n22602 = ~n3367 & ~n22406;
  assign n22603 =  a[29]  & ~n22602;
  assign n22604 = n3606 & ~n22406;
  assign n22605 = n3457 & n22402;
  assign n22606 = ~n22604 & ~n22605;
  assign n22607 = n22402 & n22406;
  assign n22608 = ~n22402 & ~n22406;
  assign n22609 = ~n22607 & ~n22608;
  assign n22610 = n3368 & ~n22609;
  assign n22611 = n22606 & ~n22610;
  assign n22612 =  a[29]  & ~n22611;
  assign n22613 =  a[29]  & ~n22612;
  assign n22614 = ~n22611 & ~n22612;
  assign n22615 = ~n22613 & ~n22614;
  assign n22616 = n22603 & ~n22615;
  assign n22617 = n3457 & n22399;
  assign n22618 = n3542 & ~n22406;
  assign n22619 = n3606 & n22402;
  assign n22620 = ~n22618 & ~n22619;
  assign n22621 = ~n22617 & n22620;
  assign n22622 = ~n3368 & n22621;
  assign n22623 = ~n22399 & n22607;
  assign n22624 = n22399 & ~n22607;
  assign n22625 = ~n22623 & ~n22624;
  assign n22626 = n22621 & n22625;
  assign n22627 = ~n22622 & ~n22626;
  assign n22628 =  a[29]  & ~n22627;
  assign n22629 = ~ a[29]  & n22627;
  assign n22630 = ~n22628 & ~n22629;
  assign n22631 = n22616 & ~n22630;
  assign n22632 = ~n7479 & ~n22406;
  assign n22633 = n22631 & ~n22632;
  assign n22634 = ~n22631 & n22632;
  assign n22635 = ~n22633 & ~n22634;
  assign n22636 = ~n22601 & ~n22635;
  assign n22637 = n22601 & n22635;
  assign n22638 = ~n22636 & ~n22637;
  assign n22639 = ~n22588 & n22638;
  assign n22640 = ~n22588 & ~n22639;
  assign n22641 = n22638 & ~n22639;
  assign n22642 = ~n22640 & ~n22641;
  assign n22643 = n3884 & n22390;
  assign n22644 = n3967 & n22396;
  assign n22645 = n4046 & n22393;
  assign n22646 = ~n22644 & ~n22645;
  assign n22647 = ~n22643 & n22646;
  assign n22648 = n22417 & ~n22419;
  assign n22649 = ~n22420 & ~n22648;
  assign n22650 = n4050 & n22649;
  assign n22651 = n22647 & ~n22650;
  assign n22652 =  a[26]  & ~n22651;
  assign n22653 = ~n22651 & ~n22652;
  assign n22654 =  a[26]  & ~n22652;
  assign n22655 = ~n22653 & ~n22654;
  assign n22656 = ~n22616 & n22630;
  assign n22657 = ~n22631 & ~n22656;
  assign n22658 = ~n22655 & n22657;
  assign n22659 = ~n22655 & ~n22658;
  assign n22660 = n22657 & ~n22658;
  assign n22661 = ~n22659 & ~n22660;
  assign n22662 = ~n22603 & n22615;
  assign n22663 = ~n22616 & ~n22662;
  assign n22664 = n3884 & n22393;
  assign n22665 = n3967 & n22399;
  assign n22666 = n4046 & n22396;
  assign n22667 = ~n22665 & ~n22666;
  assign n22668 = ~n22664 & n22667;
  assign n22669 = ~n4050 & n22668;
  assign n22670 = n22413 & ~n22415;
  assign n22671 = ~n22416 & ~n22670;
  assign n22672 = n22668 & ~n22671;
  assign n22673 = ~n22669 & ~n22672;
  assign n22674 =  a[26]  & ~n22673;
  assign n22675 = ~ a[26]  & n22673;
  assign n22676 = ~n22674 & ~n22675;
  assign n22677 = n22663 & ~n22676;
  assign n22678 = ~n3880 & ~n22406;
  assign n22679 =  a[26]  & ~n22678;
  assign n22680 = n4046 & ~n22406;
  assign n22681 = n3884 & n22402;
  assign n22682 = ~n22680 & ~n22681;
  assign n22683 = n4050 & ~n22609;
  assign n22684 = n22682 & ~n22683;
  assign n22685 =  a[26]  & ~n22684;
  assign n22686 =  a[26]  & ~n22685;
  assign n22687 = ~n22684 & ~n22685;
  assign n22688 = ~n22686 & ~n22687;
  assign n22689 = n22679 & ~n22688;
  assign n22690 = n3884 & n22399;
  assign n22691 = n3967 & ~n22406;
  assign n22692 = n4046 & n22402;
  assign n22693 = ~n22691 & ~n22692;
  assign n22694 = ~n22690 & n22693;
  assign n22695 = ~n4050 & n22694;
  assign n22696 = n22625 & n22694;
  assign n22697 = ~n22695 & ~n22696;
  assign n22698 =  a[26]  & ~n22697;
  assign n22699 = ~ a[26]  & n22697;
  assign n22700 = ~n22698 & ~n22699;
  assign n22701 = n22689 & ~n22700;
  assign n22702 = n22602 & n22701;
  assign n22703 = n22701 & ~n22702;
  assign n22704 = n22602 & ~n22702;
  assign n22705 = ~n22703 & ~n22704;
  assign n22706 = n3884 & n22396;
  assign n22707 = n3967 & n22402;
  assign n22708 = n4046 & n22399;
  assign n22709 = ~n22707 & ~n22708;
  assign n22710 = ~n22706 & n22709;
  assign n22711 = n4050 & n22595;
  assign n22712 = n22710 & ~n22711;
  assign n22713 =  a[26]  & ~n22712;
  assign n22714 =  a[26]  & ~n22713;
  assign n22715 = ~n22712 & ~n22713;
  assign n22716 = ~n22714 & ~n22715;
  assign n22717 = ~n22705 & ~n22716;
  assign n22718 = ~n22702 & ~n22717;
  assign n22719 = ~n22663 & n22676;
  assign n22720 = ~n22677 & ~n22719;
  assign n22721 = ~n22718 & n22720;
  assign n22722 = ~n22677 & ~n22721;
  assign n22723 = ~n22661 & ~n22722;
  assign n22724 = ~n22658 & ~n22723;
  assign n22725 = ~n22642 & ~n22724;
  assign n22726 = ~n22639 & ~n22725;
  assign n22727 = n3457 & n22393;
  assign n22728 = n3542 & n22399;
  assign n22729 = n3606 & n22396;
  assign n22730 = ~n22728 & ~n22729;
  assign n22731 = ~n22727 & n22730;
  assign n22732 = n3368 & n22671;
  assign n22733 = n22731 & ~n22732;
  assign n22734 =  a[29]  & ~n22733;
  assign n22735 = ~n22733 & ~n22734;
  assign n22736 =  a[29]  & ~n22734;
  assign n22737 = ~n22735 & ~n22736;
  assign n22738 = n437 & n2091;
  assign n22739 = n885 & n22738;
  assign n22740 = n108 & n22739;
  assign n22741 = n1367 & n22740;
  assign n22742 = ~n462 & n22741;
  assign n22743 = ~n149 & n22742;
  assign n22744 = ~n228 & n22743;
  assign n22745 = ~n416 & n22744;
  assign n22746 = ~n980 & n22745;
  assign n22747 = ~n791 & n22746;
  assign n22748 = ~n712 & n22747;
  assign n22749 = n3206 & n3858;
  assign n22750 = n2809 & n22749;
  assign n22751 = n4104 & n22750;
  assign n22752 = n14189 & n22751;
  assign n22753 = n804 & n22752;
  assign n22754 = n3163 & n22753;
  assign n22755 = n2276 & n22754;
  assign n22756 = n634 & n22755;
  assign n22757 = n418 & n22756;
  assign n22758 = n538 & n22757;
  assign n22759 = ~n490 & n22758;
  assign n22760 = ~n589 & n22759;
  assign n22761 = ~n163 & n22760;
  assign n22762 = ~n451 & n22761;
  assign n22763 = n735 & n2075;
  assign n22764 = n1044 & n22763;
  assign n22765 = n15956 & n22764;
  assign n22766 = n22762 & n22765;
  assign n22767 = n22748 & n22766;
  assign n22768 = n15867 & n22767;
  assign n22769 = n1161 & n22768;
  assign n22770 = n1269 & n22769;
  assign n22771 = n1180 & n22770;
  assign n22772 = n810 & n22771;
  assign n22773 = n1128 & n22772;
  assign n22774 = n341 & n22773;
  assign n22775 = ~n397 & n22774;
  assign n22776 = ~n189 & n22775;
  assign n22777 = ~n331 & n22776;
  assign n22778 = ~n144 & n22777;
  assign n22779 = ~n366 & n22778;
  assign n22780 = n3020 & n22402;
  assign n22781 = n75 & ~n22609;
  assign n22782 = n3028 & ~n22406;
  assign n22783 = ~n22781 & ~n22782;
  assign n22784 = ~n22780 & n22783;
  assign n22785 = ~n22779 & ~n22784;
  assign n22786 = ~n22779 & ~n22785;
  assign n22787 = ~n22784 & ~n22785;
  assign n22788 = ~n22786 & ~n22787;
  assign n22789 = ~n22737 & ~n22788;
  assign n22790 = ~n22737 & ~n22789;
  assign n22791 = ~n22788 & ~n22789;
  assign n22792 = ~n22790 & ~n22791;
  assign n22793 = n22631 & n22632;
  assign n22794 = ~n22636 & ~n22793;
  assign n22795 = ~n22792 & ~n22794;
  assign n22796 = ~n22792 & ~n22795;
  assign n22797 = ~n22794 & ~n22795;
  assign n22798 = ~n22796 & ~n22797;
  assign n22799 = n3884 & n22384;
  assign n22800 = n3967 & n22390;
  assign n22801 = n4046 & n22387;
  assign n22802 = ~n22800 & ~n22801;
  assign n22803 = ~n22799 & n22802;
  assign n22804 = ~n4050 & n22803;
  assign n22805 = n22425 & ~n22427;
  assign n22806 = ~n22428 & ~n22805;
  assign n22807 = n22803 & ~n22806;
  assign n22808 = ~n22804 & ~n22807;
  assign n22809 =  a[26]  & ~n22808;
  assign n22810 = ~ a[26]  & n22808;
  assign n22811 = ~n22809 & ~n22810;
  assign n22812 = ~n22798 & ~n22811;
  assign n22813 = ~n22798 & ~n22812;
  assign n22814 = ~n22811 & ~n22812;
  assign n22815 = ~n22813 & ~n22814;
  assign n22816 = ~n22726 & ~n22815;
  assign n22817 = ~n22726 & ~n22816;
  assign n22818 = ~n22815 & ~n22816;
  assign n22819 = ~n22817 & ~n22818;
  assign n22820 = ~n22575 & ~n22819;
  assign n22821 = ~n22575 & ~n22820;
  assign n22822 = ~n22819 & ~n22820;
  assign n22823 = ~n22821 & ~n22822;
  assign n22824 = n22642 & n22724;
  assign n22825 = ~n22725 & ~n22824;
  assign n22826 = n4694 & n22377;
  assign n22827 = n4533 & n22384;
  assign n22828 = n4604 & n22380;
  assign n22829 = ~n22827 & ~n22828;
  assign n22830 = ~n22826 & n22829;
  assign n22831 = ~n4536 & n22830;
  assign n22832 = ~n22433 & ~n22435;
  assign n22833 = ~n22382 & n22436;
  assign n22834 = ~n22832 & ~n22833;
  assign n22835 = n22830 & n22834;
  assign n22836 = ~n22831 & ~n22835;
  assign n22837 =  a[23]  & ~n22836;
  assign n22838 = ~ a[23]  & n22836;
  assign n22839 = ~n22837 & ~n22838;
  assign n22840 = n22825 & ~n22839;
  assign n22841 = n22661 & n22722;
  assign n22842 = ~n22723 & ~n22841;
  assign n22843 = n4694 & n22380;
  assign n22844 = n4533 & n22387;
  assign n22845 = n4604 & n22384;
  assign n22846 = ~n22844 & ~n22845;
  assign n22847 = ~n22843 & n22846;
  assign n22848 = ~n4536 & n22847;
  assign n22849 = n22429 & ~n22431;
  assign n22850 = ~n22432 & ~n22849;
  assign n22851 = n22847 & ~n22850;
  assign n22852 = ~n22848 & ~n22851;
  assign n22853 =  a[23]  & ~n22852;
  assign n22854 = ~ a[23]  & n22852;
  assign n22855 = ~n22853 & ~n22854;
  assign n22856 = n22842 & ~n22855;
  assign n22857 = n4694 & n22384;
  assign n22858 = n4533 & n22390;
  assign n22859 = n4604 & n22387;
  assign n22860 = ~n22858 & ~n22859;
  assign n22861 = ~n22857 & n22860;
  assign n22862 = n4536 & n22806;
  assign n22863 = n22861 & ~n22862;
  assign n22864 =  a[23]  & ~n22863;
  assign n22865 = ~n22863 & ~n22864;
  assign n22866 =  a[23]  & ~n22864;
  assign n22867 = ~n22865 & ~n22866;
  assign n22868 = n22718 & ~n22720;
  assign n22869 = ~n22721 & ~n22868;
  assign n22870 = ~n22867 & n22869;
  assign n22871 = ~n22867 & ~n22870;
  assign n22872 = n22869 & ~n22870;
  assign n22873 = ~n22871 & ~n22872;
  assign n22874 = ~n22705 & ~n22717;
  assign n22875 = ~n22716 & ~n22717;
  assign n22876 = ~n22874 & ~n22875;
  assign n22877 = n4694 & n22387;
  assign n22878 = n4533 & n22393;
  assign n22879 = n4604 & n22390;
  assign n22880 = ~n22878 & ~n22879;
  assign n22881 = ~n22877 & n22880;
  assign n22882 = ~n4536 & n22881;
  assign n22883 = ~n22582 & n22881;
  assign n22884 = ~n22882 & ~n22883;
  assign n22885 =  a[23]  & ~n22884;
  assign n22886 = ~ a[23]  & n22884;
  assign n22887 = ~n22885 & ~n22886;
  assign n22888 = ~n22876 & ~n22887;
  assign n22889 = n4694 & n22390;
  assign n22890 = n4533 & n22396;
  assign n22891 = n4604 & n22393;
  assign n22892 = ~n22890 & ~n22891;
  assign n22893 = ~n22889 & n22892;
  assign n22894 = n4536 & n22649;
  assign n22895 = n22893 & ~n22894;
  assign n22896 =  a[23]  & ~n22895;
  assign n22897 = ~n22895 & ~n22896;
  assign n22898 =  a[23]  & ~n22896;
  assign n22899 = ~n22897 & ~n22898;
  assign n22900 = ~n22689 & n22700;
  assign n22901 = ~n22701 & ~n22900;
  assign n22902 = ~n22899 & n22901;
  assign n22903 = ~n22899 & ~n22902;
  assign n22904 = n22901 & ~n22902;
  assign n22905 = ~n22903 & ~n22904;
  assign n22906 = ~n22679 & n22688;
  assign n22907 = ~n22689 & ~n22906;
  assign n22908 = n4694 & n22393;
  assign n22909 = n4533 & n22399;
  assign n22910 = n4604 & n22396;
  assign n22911 = ~n22909 & ~n22910;
  assign n22912 = ~n22908 & n22911;
  assign n22913 = ~n4536 & n22912;
  assign n22914 = ~n22671 & n22912;
  assign n22915 = ~n22913 & ~n22914;
  assign n22916 =  a[23]  & ~n22915;
  assign n22917 = ~ a[23]  & n22915;
  assign n22918 = ~n22916 & ~n22917;
  assign n22919 = n22907 & ~n22918;
  assign n22920 = ~n4528 & ~n22406;
  assign n22921 =  a[23]  & ~n22920;
  assign n22922 = n4604 & ~n22406;
  assign n22923 = n4694 & n22402;
  assign n22924 = ~n22922 & ~n22923;
  assign n22925 = n4536 & ~n22609;
  assign n22926 = n22924 & ~n22925;
  assign n22927 =  a[23]  & ~n22926;
  assign n22928 =  a[23]  & ~n22927;
  assign n22929 = ~n22926 & ~n22927;
  assign n22930 = ~n22928 & ~n22929;
  assign n22931 = n22921 & ~n22930;
  assign n22932 = n4694 & n22399;
  assign n22933 = n4533 & ~n22406;
  assign n22934 = n4604 & n22402;
  assign n22935 = ~n22933 & ~n22934;
  assign n22936 = ~n22932 & n22935;
  assign n22937 = ~n4536 & n22936;
  assign n22938 = n22625 & n22936;
  assign n22939 = ~n22937 & ~n22938;
  assign n22940 =  a[23]  & ~n22939;
  assign n22941 = ~ a[23]  & n22939;
  assign n22942 = ~n22940 & ~n22941;
  assign n22943 = n22931 & ~n22942;
  assign n22944 = n22678 & n22943;
  assign n22945 = n22943 & ~n22944;
  assign n22946 = n22678 & ~n22944;
  assign n22947 = ~n22945 & ~n22946;
  assign n22948 = n4694 & n22396;
  assign n22949 = n4533 & n22402;
  assign n22950 = n4604 & n22399;
  assign n22951 = ~n22949 & ~n22950;
  assign n22952 = ~n22948 & n22951;
  assign n22953 = n4536 & n22595;
  assign n22954 = n22952 & ~n22953;
  assign n22955 =  a[23]  & ~n22954;
  assign n22956 =  a[23]  & ~n22955;
  assign n22957 = ~n22954 & ~n22955;
  assign n22958 = ~n22956 & ~n22957;
  assign n22959 = ~n22947 & ~n22958;
  assign n22960 = ~n22944 & ~n22959;
  assign n22961 = ~n22907 & n22918;
  assign n22962 = ~n22919 & ~n22961;
  assign n22963 = ~n22960 & n22962;
  assign n22964 = ~n22919 & ~n22963;
  assign n22965 = ~n22905 & ~n22964;
  assign n22966 = ~n22902 & ~n22965;
  assign n22967 = n22876 & n22887;
  assign n22968 = ~n22888 & ~n22967;
  assign n22969 = ~n22966 & n22968;
  assign n22970 = ~n22888 & ~n22969;
  assign n22971 = ~n22873 & ~n22970;
  assign n22972 = ~n22870 & ~n22971;
  assign n22973 = n22842 & ~n22856;
  assign n22974 = ~n22855 & ~n22856;
  assign n22975 = ~n22973 & ~n22974;
  assign n22976 = ~n22972 & ~n22975;
  assign n22977 = ~n22856 & ~n22976;
  assign n22978 = ~n22825 & n22839;
  assign n22979 = ~n22840 & ~n22978;
  assign n22980 = ~n22977 & n22979;
  assign n22981 = ~n22840 & ~n22980;
  assign n22982 = n22823 & n22981;
  assign n22983 = ~n22823 & ~n22981;
  assign n22984 = ~n22982 & ~n22983;
  assign n22985 = n5496 & n22365;
  assign n22986 = n4935 & n22371;
  assign n22987 = n5407 & n22368;
  assign n22988 = ~n22986 & ~n22987;
  assign n22989 = ~n22985 & n22988;
  assign n22990 = ~n4938 & n22989;
  assign n22991 = ~n22448 & ~n22451;
  assign n22992 = ~n22449 & n22452;
  assign n22993 = ~n22991 & ~n22992;
  assign n22994 = n22989 & n22993;
  assign n22995 = ~n22990 & ~n22994;
  assign n22996 =  a[20]  & ~n22995;
  assign n22997 = ~ a[20]  & n22995;
  assign n22998 = ~n22996 & ~n22997;
  assign n22999 = n22984 & ~n22998;
  assign n23000 = n5496 & n22368;
  assign n23001 = n4935 & n22374;
  assign n23002 = n5407 & n22371;
  assign n23003 = ~n23001 & ~n23002;
  assign n23004 = ~n23000 & n23003;
  assign n23005 = n22444 & ~n22446;
  assign n23006 = ~n22447 & ~n23005;
  assign n23007 = n4938 & n23006;
  assign n23008 = n23004 & ~n23007;
  assign n23009 =  a[20]  & ~n23008;
  assign n23010 = ~n23008 & ~n23009;
  assign n23011 =  a[20]  & ~n23009;
  assign n23012 = ~n23010 & ~n23011;
  assign n23013 = n22977 & ~n22979;
  assign n23014 = ~n22980 & ~n23013;
  assign n23015 = ~n23012 & n23014;
  assign n23016 = ~n23012 & ~n23015;
  assign n23017 = n23014 & ~n23015;
  assign n23018 = ~n23016 & ~n23017;
  assign n23019 = n5496 & n22371;
  assign n23020 = n4935 & n22377;
  assign n23021 = n5407 & n22374;
  assign n23022 = ~n23020 & ~n23021;
  assign n23023 = ~n23019 & n23022;
  assign n23024 = n22440 & ~n22442;
  assign n23025 = ~n22443 & ~n23024;
  assign n23026 = n4938 & n23025;
  assign n23027 = n23023 & ~n23026;
  assign n23028 =  a[20]  & ~n23027;
  assign n23029 = ~n23027 & ~n23028;
  assign n23030 =  a[20]  & ~n23028;
  assign n23031 = ~n23029 & ~n23030;
  assign n23032 = ~n22972 & ~n22976;
  assign n23033 = ~n22975 & ~n22976;
  assign n23034 = ~n23032 & ~n23033;
  assign n23035 = ~n23031 & ~n23034;
  assign n23036 = ~n23031 & ~n23035;
  assign n23037 = ~n23034 & ~n23035;
  assign n23038 = ~n23036 & ~n23037;
  assign n23039 = n22873 & n22970;
  assign n23040 = ~n22971 & ~n23039;
  assign n23041 = n5496 & n22374;
  assign n23042 = n4935 & n22380;
  assign n23043 = n5407 & n22377;
  assign n23044 = ~n23042 & ~n23043;
  assign n23045 = ~n23041 & n23044;
  assign n23046 = ~n4938 & n23045;
  assign n23047 = ~n22569 & n23045;
  assign n23048 = ~n23046 & ~n23047;
  assign n23049 =  a[20]  & ~n23048;
  assign n23050 = ~ a[20]  & n23048;
  assign n23051 = ~n23049 & ~n23050;
  assign n23052 = n23040 & ~n23051;
  assign n23053 = n22966 & ~n22968;
  assign n23054 = ~n22969 & ~n23053;
  assign n23055 = n5496 & n22377;
  assign n23056 = n4935 & n22384;
  assign n23057 = n5407 & n22380;
  assign n23058 = ~n23056 & ~n23057;
  assign n23059 = ~n23055 & n23058;
  assign n23060 = ~n4938 & n23059;
  assign n23061 = n22834 & n23059;
  assign n23062 = ~n23060 & ~n23061;
  assign n23063 =  a[20]  & ~n23062;
  assign n23064 = ~ a[20]  & n23062;
  assign n23065 = ~n23063 & ~n23064;
  assign n23066 = n23054 & ~n23065;
  assign n23067 = n22905 & n22964;
  assign n23068 = ~n22965 & ~n23067;
  assign n23069 = n5496 & n22380;
  assign n23070 = n4935 & n22387;
  assign n23071 = n5407 & n22384;
  assign n23072 = ~n23070 & ~n23071;
  assign n23073 = ~n23069 & n23072;
  assign n23074 = ~n4938 & n23073;
  assign n23075 = ~n22850 & n23073;
  assign n23076 = ~n23074 & ~n23075;
  assign n23077 =  a[20]  & ~n23076;
  assign n23078 = ~ a[20]  & n23076;
  assign n23079 = ~n23077 & ~n23078;
  assign n23080 = n23068 & ~n23079;
  assign n23081 = n5496 & n22384;
  assign n23082 = n4935 & n22390;
  assign n23083 = n5407 & n22387;
  assign n23084 = ~n23082 & ~n23083;
  assign n23085 = ~n23081 & n23084;
  assign n23086 = n4938 & n22806;
  assign n23087 = n23085 & ~n23086;
  assign n23088 =  a[20]  & ~n23087;
  assign n23089 = ~n23087 & ~n23088;
  assign n23090 =  a[20]  & ~n23088;
  assign n23091 = ~n23089 & ~n23090;
  assign n23092 = n22960 & ~n22962;
  assign n23093 = ~n22963 & ~n23092;
  assign n23094 = ~n23091 & n23093;
  assign n23095 = ~n23091 & ~n23094;
  assign n23096 = n23093 & ~n23094;
  assign n23097 = ~n23095 & ~n23096;
  assign n23098 = ~n22947 & ~n22959;
  assign n23099 = ~n22958 & ~n22959;
  assign n23100 = ~n23098 & ~n23099;
  assign n23101 = n5496 & n22387;
  assign n23102 = n4935 & n22393;
  assign n23103 = n5407 & n22390;
  assign n23104 = ~n23102 & ~n23103;
  assign n23105 = ~n23101 & n23104;
  assign n23106 = ~n4938 & n23105;
  assign n23107 = ~n22582 & n23105;
  assign n23108 = ~n23106 & ~n23107;
  assign n23109 =  a[20]  & ~n23108;
  assign n23110 = ~ a[20]  & n23108;
  assign n23111 = ~n23109 & ~n23110;
  assign n23112 = ~n23100 & ~n23111;
  assign n23113 = n5496 & n22390;
  assign n23114 = n4935 & n22396;
  assign n23115 = n5407 & n22393;
  assign n23116 = ~n23114 & ~n23115;
  assign n23117 = ~n23113 & n23116;
  assign n23118 = n4938 & n22649;
  assign n23119 = n23117 & ~n23118;
  assign n23120 =  a[20]  & ~n23119;
  assign n23121 = ~n23119 & ~n23120;
  assign n23122 =  a[20]  & ~n23120;
  assign n23123 = ~n23121 & ~n23122;
  assign n23124 = ~n22931 & n22942;
  assign n23125 = ~n22943 & ~n23124;
  assign n23126 = ~n23123 & n23125;
  assign n23127 = ~n23123 & ~n23126;
  assign n23128 = n23125 & ~n23126;
  assign n23129 = ~n23127 & ~n23128;
  assign n23130 = ~n22921 & n22930;
  assign n23131 = ~n22931 & ~n23130;
  assign n23132 = n5496 & n22393;
  assign n23133 = n4935 & n22399;
  assign n23134 = n5407 & n22396;
  assign n23135 = ~n23133 & ~n23134;
  assign n23136 = ~n23132 & n23135;
  assign n23137 = ~n4938 & n23136;
  assign n23138 = ~n22671 & n23136;
  assign n23139 = ~n23137 & ~n23138;
  assign n23140 =  a[20]  & ~n23139;
  assign n23141 = ~ a[20]  & n23139;
  assign n23142 = ~n23140 & ~n23141;
  assign n23143 = n23131 & ~n23142;
  assign n23144 = n5407 & ~n22406;
  assign n23145 = n5496 & n22402;
  assign n23146 = ~n23144 & ~n23145;
  assign n23147 = n4938 & ~n22609;
  assign n23148 = n23146 & ~n23147;
  assign n23149 =  a[20]  & ~n23148;
  assign n23150 =  a[20]  & ~n23149;
  assign n23151 = ~n23148 & ~n23149;
  assign n23152 = ~n23150 & ~n23151;
  assign n23153 = ~n4933 & ~n22406;
  assign n23154 =  a[20]  & ~n23153;
  assign n23155 = ~n23152 & n23154;
  assign n23156 = n5496 & n22399;
  assign n23157 = n4935 & ~n22406;
  assign n23158 = n5407 & n22402;
  assign n23159 = ~n23157 & ~n23158;
  assign n23160 = ~n23156 & n23159;
  assign n23161 = ~n4938 & n23160;
  assign n23162 = n22625 & n23160;
  assign n23163 = ~n23161 & ~n23162;
  assign n23164 =  a[20]  & ~n23163;
  assign n23165 = ~ a[20]  & n23163;
  assign n23166 = ~n23164 & ~n23165;
  assign n23167 = n23155 & ~n23166;
  assign n23168 = n22920 & n23167;
  assign n23169 = n23167 & ~n23168;
  assign n23170 = n22920 & ~n23168;
  assign n23171 = ~n23169 & ~n23170;
  assign n23172 = n5496 & n22396;
  assign n23173 = n4935 & n22402;
  assign n23174 = n5407 & n22399;
  assign n23175 = ~n23173 & ~n23174;
  assign n23176 = ~n23172 & n23175;
  assign n23177 = n4938 & n22595;
  assign n23178 = n23176 & ~n23177;
  assign n23179 =  a[20]  & ~n23178;
  assign n23180 =  a[20]  & ~n23179;
  assign n23181 = ~n23178 & ~n23179;
  assign n23182 = ~n23180 & ~n23181;
  assign n23183 = ~n23171 & ~n23182;
  assign n23184 = ~n23168 & ~n23183;
  assign n23185 = ~n23131 & n23142;
  assign n23186 = ~n23143 & ~n23185;
  assign n23187 = ~n23184 & n23186;
  assign n23188 = ~n23143 & ~n23187;
  assign n23189 = ~n23129 & ~n23188;
  assign n23190 = ~n23126 & ~n23189;
  assign n23191 = n23100 & n23111;
  assign n23192 = ~n23112 & ~n23191;
  assign n23193 = ~n23190 & n23192;
  assign n23194 = ~n23112 & ~n23193;
  assign n23195 = ~n23097 & ~n23194;
  assign n23196 = ~n23094 & ~n23195;
  assign n23197 = n23068 & ~n23080;
  assign n23198 = ~n23079 & ~n23080;
  assign n23199 = ~n23197 & ~n23198;
  assign n23200 = ~n23196 & ~n23199;
  assign n23201 = ~n23080 & ~n23200;
  assign n23202 = n23054 & ~n23066;
  assign n23203 = ~n23065 & ~n23066;
  assign n23204 = ~n23202 & ~n23203;
  assign n23205 = ~n23201 & ~n23204;
  assign n23206 = ~n23066 & ~n23205;
  assign n23207 = ~n23040 & n23051;
  assign n23208 = ~n23052 & ~n23207;
  assign n23209 = ~n23206 & n23208;
  assign n23210 = ~n23052 & ~n23209;
  assign n23211 = ~n23038 & ~n23210;
  assign n23212 = ~n23035 & ~n23211;
  assign n23213 = ~n23018 & ~n23212;
  assign n23214 = ~n23015 & ~n23213;
  assign n23215 = n22984 & ~n22999;
  assign n23216 = ~n22998 & ~n22999;
  assign n23217 = ~n23215 & ~n23216;
  assign n23218 = ~n23214 & ~n23217;
  assign n23219 = ~n22999 & ~n23218;
  assign n23220 = n4694 & n22371;
  assign n23221 = n4533 & n22377;
  assign n23222 = n4604 & n22374;
  assign n23223 = ~n23221 & ~n23222;
  assign n23224 = ~n23220 & n23223;
  assign n23225 = n4536 & n23025;
  assign n23226 = n23224 & ~n23225;
  assign n23227 =  a[23]  & ~n23226;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 =  a[23]  & ~n23227;
  assign n23230 = ~n23228 & ~n23229;
  assign n23231 = ~n22812 & ~n22816;
  assign n23232 = n3457 & n22390;
  assign n23233 = n3542 & n22396;
  assign n23234 = n3606 & n22393;
  assign n23235 = ~n23233 & ~n23234;
  assign n23236 = ~n23232 & n23235;
  assign n23237 = n3368 & n22649;
  assign n23238 = n23236 & ~n23237;
  assign n23239 =  a[29]  & ~n23238;
  assign n23240 = ~n23238 & ~n23239;
  assign n23241 =  a[29]  & ~n23239;
  assign n23242 = ~n23240 & ~n23241;
  assign n23243 = n75 & ~n22625;
  assign n23244 = n3020 & n22399;
  assign n23245 = n3023 & ~n22406;
  assign n23246 = n3028 & n22402;
  assign n23247 = ~n23245 & ~n23246;
  assign n23248 = ~n23244 & n23247;
  assign n23249 = ~n23243 & n23248;
  assign n23250 = ~n233 & ~n332;
  assign n23251 = ~n86 & n23250;
  assign n23252 = n13774 & n23251;
  assign n23253 = n3041 & n23252;
  assign n23254 = n12387 & n23253;
  assign n23255 = n732 & n23254;
  assign n23256 = n3261 & n23255;
  assign n23257 = n6625 & n23256;
  assign n23258 = n5209 & n23257;
  assign n23259 = n967 & n23258;
  assign n23260 = n294 & n23259;
  assign n23261 = n1129 & n23260;
  assign n23262 = n731 & n23261;
  assign n23263 = n15867 & n23262;
  assign n23264 = ~n420 & n23263;
  assign n23265 = ~n280 & n23264;
  assign n23266 = ~n228 & n23265;
  assign n23267 = ~n980 & n23266;
  assign n23268 = ~n673 & n23267;
  assign n23269 = ~n567 & n23268;
  assign n23270 = n22785 & ~n23269;
  assign n23271 = ~n22785 & n23269;
  assign n23272 = ~n23270 & ~n23271;
  assign n23273 = ~n23249 & n23272;
  assign n23274 = ~n23249 & ~n23273;
  assign n23275 = n23272 & ~n23273;
  assign n23276 = ~n23274 & ~n23275;
  assign n23277 = ~n23242 & ~n23276;
  assign n23278 = ~n23242 & ~n23277;
  assign n23279 = ~n23276 & ~n23277;
  assign n23280 = ~n23278 & ~n23279;
  assign n23281 = ~n22789 & ~n22795;
  assign n23282 = n23280 & n23281;
  assign n23283 = ~n23280 & ~n23281;
  assign n23284 = ~n23282 & ~n23283;
  assign n23285 = n3884 & n22380;
  assign n23286 = n3967 & n22387;
  assign n23287 = n4046 & n22384;
  assign n23288 = ~n23286 & ~n23287;
  assign n23289 = ~n23285 & n23288;
  assign n23290 = ~n4050 & n23289;
  assign n23291 = ~n22850 & n23289;
  assign n23292 = ~n23290 & ~n23291;
  assign n23293 =  a[26]  & ~n23292;
  assign n23294 = ~ a[26]  & n23292;
  assign n23295 = ~n23293 & ~n23294;
  assign n23296 = n23284 & ~n23295;
  assign n23297 = n23284 & ~n23296;
  assign n23298 = ~n23295 & ~n23296;
  assign n23299 = ~n23297 & ~n23298;
  assign n23300 = ~n23231 & ~n23299;
  assign n23301 = ~n23231 & ~n23300;
  assign n23302 = ~n23299 & ~n23300;
  assign n23303 = ~n23301 & ~n23302;
  assign n23304 = ~n23230 & ~n23303;
  assign n23305 = ~n23230 & ~n23304;
  assign n23306 = ~n23303 & ~n23304;
  assign n23307 = ~n23305 & ~n23306;
  assign n23308 = ~n22820 & ~n22983;
  assign n23309 = n23307 & n23308;
  assign n23310 = ~n23307 & ~n23308;
  assign n23311 = ~n23309 & ~n23310;
  assign n23312 = n5496 & n22362;
  assign n23313 = n4935 & n22368;
  assign n23314 = n5407 & n22365;
  assign n23315 = ~n23313 & ~n23314;
  assign n23316 = ~n23312 & n23315;
  assign n23317 = ~n4938 & n23316;
  assign n23318 = ~n22452 & ~n22455;
  assign n23319 = ~n22453 & n22456;
  assign n23320 = ~n23318 & ~n23319;
  assign n23321 = n23316 & n23320;
  assign n23322 = ~n23317 & ~n23321;
  assign n23323 =  a[20]  & ~n23322;
  assign n23324 = ~ a[20]  & n23322;
  assign n23325 = ~n23323 & ~n23324;
  assign n23326 = n23311 & ~n23325;
  assign n23327 = n23311 & ~n23326;
  assign n23328 = ~n23325 & ~n23326;
  assign n23329 = ~n23327 & ~n23328;
  assign n23330 = ~n23219 & ~n23329;
  assign n23331 = ~n23219 & ~n23330;
  assign n23332 = ~n23329 & ~n23330;
  assign n23333 = ~n23331 & ~n23332;
  assign n23334 = ~n22562 & ~n23333;
  assign n23335 = ~n22562 & ~n23334;
  assign n23336 = ~n23333 & ~n23334;
  assign n23337 = ~n23335 & ~n23336;
  assign n23338 = n6233 & n22356;
  assign n23339 = n5663 & n22362;
  assign n23340 = n5939 & n22359;
  assign n23341 = ~n23339 & ~n23340;
  assign n23342 = ~n23338 & n23341;
  assign n23343 = ~n22460 & ~n22463;
  assign n23344 = ~n22461 & n22464;
  assign n23345 = ~n23343 & ~n23344;
  assign n23346 = n5666 & ~n23345;
  assign n23347 = n23342 & ~n23346;
  assign n23348 =  a[17]  & ~n23347;
  assign n23349 = ~n23347 & ~n23348;
  assign n23350 =  a[17]  & ~n23348;
  assign n23351 = ~n23349 & ~n23350;
  assign n23352 = ~n23214 & ~n23218;
  assign n23353 = ~n23217 & ~n23218;
  assign n23354 = ~n23352 & ~n23353;
  assign n23355 = ~n23351 & ~n23354;
  assign n23356 = ~n23351 & ~n23355;
  assign n23357 = ~n23354 & ~n23355;
  assign n23358 = ~n23356 & ~n23357;
  assign n23359 = n23018 & n23212;
  assign n23360 = ~n23213 & ~n23359;
  assign n23361 = n6233 & n22359;
  assign n23362 = n5663 & n22365;
  assign n23363 = n5939 & n22362;
  assign n23364 = ~n23362 & ~n23363;
  assign n23365 = ~n23361 & n23364;
  assign n23366 = ~n5666 & n23365;
  assign n23367 = n22456 & ~n22458;
  assign n23368 = ~n22459 & ~n23367;
  assign n23369 = n23365 & ~n23368;
  assign n23370 = ~n23366 & ~n23369;
  assign n23371 =  a[17]  & ~n23370;
  assign n23372 = ~ a[17]  & n23370;
  assign n23373 = ~n23371 & ~n23372;
  assign n23374 = n23360 & ~n23373;
  assign n23375 = n23038 & n23210;
  assign n23376 = ~n23211 & ~n23375;
  assign n23377 = n6233 & n22362;
  assign n23378 = n5663 & n22368;
  assign n23379 = n5939 & n22365;
  assign n23380 = ~n23378 & ~n23379;
  assign n23381 = ~n23377 & n23380;
  assign n23382 = ~n5666 & n23381;
  assign n23383 = n23320 & n23381;
  assign n23384 = ~n23382 & ~n23383;
  assign n23385 =  a[17]  & ~n23384;
  assign n23386 = ~ a[17]  & n23384;
  assign n23387 = ~n23385 & ~n23386;
  assign n23388 = n23376 & ~n23387;
  assign n23389 = n6233 & n22365;
  assign n23390 = n5663 & n22371;
  assign n23391 = n5939 & n22368;
  assign n23392 = ~n23390 & ~n23391;
  assign n23393 = ~n23389 & n23392;
  assign n23394 = n5666 & ~n22993;
  assign n23395 = n23393 & ~n23394;
  assign n23396 =  a[17]  & ~n23395;
  assign n23397 = ~n23395 & ~n23396;
  assign n23398 =  a[17]  & ~n23396;
  assign n23399 = ~n23397 & ~n23398;
  assign n23400 = n23206 & ~n23208;
  assign n23401 = ~n23209 & ~n23400;
  assign n23402 = ~n23399 & n23401;
  assign n23403 = ~n23399 & ~n23402;
  assign n23404 = n23401 & ~n23402;
  assign n23405 = ~n23403 & ~n23404;
  assign n23406 = n6233 & n22368;
  assign n23407 = n5663 & n22374;
  assign n23408 = n5939 & n22371;
  assign n23409 = ~n23407 & ~n23408;
  assign n23410 = ~n23406 & n23409;
  assign n23411 = n5666 & n23006;
  assign n23412 = n23410 & ~n23411;
  assign n23413 =  a[17]  & ~n23412;
  assign n23414 = ~n23412 & ~n23413;
  assign n23415 =  a[17]  & ~n23413;
  assign n23416 = ~n23414 & ~n23415;
  assign n23417 = ~n23201 & ~n23205;
  assign n23418 = ~n23204 & ~n23205;
  assign n23419 = ~n23417 & ~n23418;
  assign n23420 = ~n23416 & ~n23419;
  assign n23421 = ~n23416 & ~n23420;
  assign n23422 = ~n23419 & ~n23420;
  assign n23423 = ~n23421 & ~n23422;
  assign n23424 = n6233 & n22371;
  assign n23425 = n5663 & n22377;
  assign n23426 = n5939 & n22374;
  assign n23427 = ~n23425 & ~n23426;
  assign n23428 = ~n23424 & n23427;
  assign n23429 = n5666 & n23025;
  assign n23430 = n23428 & ~n23429;
  assign n23431 =  a[17]  & ~n23430;
  assign n23432 = ~n23430 & ~n23431;
  assign n23433 =  a[17]  & ~n23431;
  assign n23434 = ~n23432 & ~n23433;
  assign n23435 = ~n23196 & ~n23200;
  assign n23436 = ~n23199 & ~n23200;
  assign n23437 = ~n23435 & ~n23436;
  assign n23438 = ~n23434 & ~n23437;
  assign n23439 = ~n23434 & ~n23438;
  assign n23440 = ~n23437 & ~n23438;
  assign n23441 = ~n23439 & ~n23440;
  assign n23442 = n23097 & n23194;
  assign n23443 = ~n23195 & ~n23442;
  assign n23444 = n6233 & n22374;
  assign n23445 = n5663 & n22380;
  assign n23446 = n5939 & n22377;
  assign n23447 = ~n23445 & ~n23446;
  assign n23448 = ~n23444 & n23447;
  assign n23449 = ~n5666 & n23448;
  assign n23450 = ~n22569 & n23448;
  assign n23451 = ~n23449 & ~n23450;
  assign n23452 =  a[17]  & ~n23451;
  assign n23453 = ~ a[17]  & n23451;
  assign n23454 = ~n23452 & ~n23453;
  assign n23455 = n23443 & ~n23454;
  assign n23456 = n23190 & ~n23192;
  assign n23457 = ~n23193 & ~n23456;
  assign n23458 = n6233 & n22377;
  assign n23459 = n5663 & n22384;
  assign n23460 = n5939 & n22380;
  assign n23461 = ~n23459 & ~n23460;
  assign n23462 = ~n23458 & n23461;
  assign n23463 = ~n5666 & n23462;
  assign n23464 = n22834 & n23462;
  assign n23465 = ~n23463 & ~n23464;
  assign n23466 =  a[17]  & ~n23465;
  assign n23467 = ~ a[17]  & n23465;
  assign n23468 = ~n23466 & ~n23467;
  assign n23469 = n23457 & ~n23468;
  assign n23470 = n23129 & n23188;
  assign n23471 = ~n23189 & ~n23470;
  assign n23472 = n6233 & n22380;
  assign n23473 = n5663 & n22387;
  assign n23474 = n5939 & n22384;
  assign n23475 = ~n23473 & ~n23474;
  assign n23476 = ~n23472 & n23475;
  assign n23477 = ~n5666 & n23476;
  assign n23478 = ~n22850 & n23476;
  assign n23479 = ~n23477 & ~n23478;
  assign n23480 =  a[17]  & ~n23479;
  assign n23481 = ~ a[17]  & n23479;
  assign n23482 = ~n23480 & ~n23481;
  assign n23483 = n23471 & ~n23482;
  assign n23484 = n6233 & n22384;
  assign n23485 = n5663 & n22390;
  assign n23486 = n5939 & n22387;
  assign n23487 = ~n23485 & ~n23486;
  assign n23488 = ~n23484 & n23487;
  assign n23489 = n5666 & n22806;
  assign n23490 = n23488 & ~n23489;
  assign n23491 =  a[17]  & ~n23490;
  assign n23492 = ~n23490 & ~n23491;
  assign n23493 =  a[17]  & ~n23491;
  assign n23494 = ~n23492 & ~n23493;
  assign n23495 = n23184 & ~n23186;
  assign n23496 = ~n23187 & ~n23495;
  assign n23497 = ~n23494 & n23496;
  assign n23498 = ~n23494 & ~n23497;
  assign n23499 = n23496 & ~n23497;
  assign n23500 = ~n23498 & ~n23499;
  assign n23501 = ~n23171 & ~n23183;
  assign n23502 = ~n23182 & ~n23183;
  assign n23503 = ~n23501 & ~n23502;
  assign n23504 = n6233 & n22387;
  assign n23505 = n5663 & n22393;
  assign n23506 = n5939 & n22390;
  assign n23507 = ~n23505 & ~n23506;
  assign n23508 = ~n23504 & n23507;
  assign n23509 = ~n5666 & n23508;
  assign n23510 = ~n22582 & n23508;
  assign n23511 = ~n23509 & ~n23510;
  assign n23512 =  a[17]  & ~n23511;
  assign n23513 = ~ a[17]  & n23511;
  assign n23514 = ~n23512 & ~n23513;
  assign n23515 = ~n23503 & ~n23514;
  assign n23516 = n6233 & n22390;
  assign n23517 = n5663 & n22396;
  assign n23518 = n5939 & n22393;
  assign n23519 = ~n23517 & ~n23518;
  assign n23520 = ~n23516 & n23519;
  assign n23521 = n5666 & n22649;
  assign n23522 = n23520 & ~n23521;
  assign n23523 =  a[17]  & ~n23522;
  assign n23524 = ~n23522 & ~n23523;
  assign n23525 =  a[17]  & ~n23523;
  assign n23526 = ~n23524 & ~n23525;
  assign n23527 = ~n23155 & n23166;
  assign n23528 = ~n23167 & ~n23527;
  assign n23529 = ~n23526 & n23528;
  assign n23530 = ~n23526 & ~n23529;
  assign n23531 = n23528 & ~n23529;
  assign n23532 = ~n23530 & ~n23531;
  assign n23533 = n23152 & ~n23154;
  assign n23534 = ~n23155 & ~n23533;
  assign n23535 = n6233 & n22393;
  assign n23536 = n5663 & n22399;
  assign n23537 = n5939 & n22396;
  assign n23538 = ~n23536 & ~n23537;
  assign n23539 = ~n23535 & n23538;
  assign n23540 = ~n5666 & n23539;
  assign n23541 = ~n22671 & n23539;
  assign n23542 = ~n23540 & ~n23541;
  assign n23543 =  a[17]  & ~n23542;
  assign n23544 = ~ a[17]  & n23542;
  assign n23545 = ~n23543 & ~n23544;
  assign n23546 = n23534 & ~n23545;
  assign n23547 = n5939 & ~n22406;
  assign n23548 = n6233 & n22402;
  assign n23549 = ~n23547 & ~n23548;
  assign n23550 = n5666 & ~n22609;
  assign n23551 = n23549 & ~n23550;
  assign n23552 =  a[17]  & ~n23551;
  assign n23553 =  a[17]  & ~n23552;
  assign n23554 = ~n23551 & ~n23552;
  assign n23555 = ~n23553 & ~n23554;
  assign n23556 = ~n5658 & ~n22406;
  assign n23557 =  a[17]  & ~n23556;
  assign n23558 = ~n23555 & n23557;
  assign n23559 = n6233 & n22399;
  assign n23560 = n5663 & ~n22406;
  assign n23561 = n5939 & n22402;
  assign n23562 = ~n23560 & ~n23561;
  assign n23563 = ~n23559 & n23562;
  assign n23564 = ~n5666 & n23563;
  assign n23565 = n22625 & n23563;
  assign n23566 = ~n23564 & ~n23565;
  assign n23567 =  a[17]  & ~n23566;
  assign n23568 = ~ a[17]  & n23566;
  assign n23569 = ~n23567 & ~n23568;
  assign n23570 = n23558 & ~n23569;
  assign n23571 = n23153 & n23570;
  assign n23572 = n23570 & ~n23571;
  assign n23573 = n23153 & ~n23571;
  assign n23574 = ~n23572 & ~n23573;
  assign n23575 = n6233 & n22396;
  assign n23576 = n5663 & n22402;
  assign n23577 = n5939 & n22399;
  assign n23578 = ~n23576 & ~n23577;
  assign n23579 = ~n23575 & n23578;
  assign n23580 = n5666 & n22595;
  assign n23581 = n23579 & ~n23580;
  assign n23582 =  a[17]  & ~n23581;
  assign n23583 =  a[17]  & ~n23582;
  assign n23584 = ~n23581 & ~n23582;
  assign n23585 = ~n23583 & ~n23584;
  assign n23586 = ~n23574 & ~n23585;
  assign n23587 = ~n23571 & ~n23586;
  assign n23588 = ~n23534 & n23545;
  assign n23589 = ~n23546 & ~n23588;
  assign n23590 = ~n23587 & n23589;
  assign n23591 = ~n23546 & ~n23590;
  assign n23592 = ~n23532 & ~n23591;
  assign n23593 = ~n23529 & ~n23592;
  assign n23594 = n23503 & n23514;
  assign n23595 = ~n23515 & ~n23594;
  assign n23596 = ~n23593 & n23595;
  assign n23597 = ~n23515 & ~n23596;
  assign n23598 = ~n23500 & ~n23597;
  assign n23599 = ~n23497 & ~n23598;
  assign n23600 = n23471 & ~n23483;
  assign n23601 = ~n23482 & ~n23483;
  assign n23602 = ~n23600 & ~n23601;
  assign n23603 = ~n23599 & ~n23602;
  assign n23604 = ~n23483 & ~n23603;
  assign n23605 = n23457 & ~n23469;
  assign n23606 = ~n23468 & ~n23469;
  assign n23607 = ~n23605 & ~n23606;
  assign n23608 = ~n23604 & ~n23607;
  assign n23609 = ~n23469 & ~n23608;
  assign n23610 = ~n23443 & n23454;
  assign n23611 = ~n23455 & ~n23610;
  assign n23612 = ~n23609 & n23611;
  assign n23613 = ~n23455 & ~n23612;
  assign n23614 = ~n23441 & ~n23613;
  assign n23615 = ~n23438 & ~n23614;
  assign n23616 = ~n23423 & ~n23615;
  assign n23617 = ~n23420 & ~n23616;
  assign n23618 = ~n23405 & ~n23617;
  assign n23619 = ~n23402 & ~n23618;
  assign n23620 = n23376 & ~n23388;
  assign n23621 = ~n23387 & ~n23388;
  assign n23622 = ~n23620 & ~n23621;
  assign n23623 = ~n23619 & ~n23622;
  assign n23624 = ~n23388 & ~n23623;
  assign n23625 = ~n23360 & n23373;
  assign n23626 = ~n23374 & ~n23625;
  assign n23627 = ~n23624 & n23626;
  assign n23628 = ~n23374 & ~n23627;
  assign n23629 = ~n23358 & ~n23628;
  assign n23630 = ~n23355 & ~n23629;
  assign n23631 = n23337 & n23630;
  assign n23632 = ~n23337 & ~n23630;
  assign n23633 = ~n23631 & ~n23632;
  assign n23634 = n7101 & n22344;
  assign n23635 = n6402 & n22350;
  assign n23636 = n6951 & n22347;
  assign n23637 = ~n23635 & ~n23636;
  assign n23638 = ~n23634 & n23637;
  assign n23639 = ~n6397 & n23638;
  assign n23640 = ~n22476 & ~n22479;
  assign n23641 = ~n22477 & n22480;
  assign n23642 = ~n23640 & ~n23641;
  assign n23643 = n23638 & n23642;
  assign n23644 = ~n23639 & ~n23643;
  assign n23645 =  a[14]  & ~n23644;
  assign n23646 = ~ a[14]  & n23644;
  assign n23647 = ~n23645 & ~n23646;
  assign n23648 = n23633 & ~n23647;
  assign n23649 = n23358 & n23628;
  assign n23650 = ~n23629 & ~n23649;
  assign n23651 = n7101 & n22347;
  assign n23652 = n6402 & n22353;
  assign n23653 = n6951 & n22350;
  assign n23654 = ~n23652 & ~n23653;
  assign n23655 = ~n23651 & n23654;
  assign n23656 = ~n6397 & n23655;
  assign n23657 = ~n22472 & ~n22475;
  assign n23658 = ~n22473 & n22476;
  assign n23659 = ~n23657 & ~n23658;
  assign n23660 = n23655 & n23659;
  assign n23661 = ~n23656 & ~n23660;
  assign n23662 =  a[14]  & ~n23661;
  assign n23663 = ~ a[14]  & n23661;
  assign n23664 = ~n23662 & ~n23663;
  assign n23665 = n23650 & ~n23664;
  assign n23666 = n7101 & n22350;
  assign n23667 = n6402 & n22356;
  assign n23668 = n6951 & n22353;
  assign n23669 = ~n23667 & ~n23668;
  assign n23670 = ~n23666 & n23669;
  assign n23671 = n22468 & ~n22470;
  assign n23672 = ~n22471 & ~n23671;
  assign n23673 = n6397 & n23672;
  assign n23674 = n23670 & ~n23673;
  assign n23675 =  a[14]  & ~n23674;
  assign n23676 = ~n23674 & ~n23675;
  assign n23677 =  a[14]  & ~n23675;
  assign n23678 = ~n23676 & ~n23677;
  assign n23679 = n23624 & ~n23626;
  assign n23680 = ~n23627 & ~n23679;
  assign n23681 = ~n23678 & n23680;
  assign n23682 = ~n23678 & ~n23681;
  assign n23683 = n23680 & ~n23681;
  assign n23684 = ~n23682 & ~n23683;
  assign n23685 = n7101 & n22353;
  assign n23686 = n6402 & n22359;
  assign n23687 = n6951 & n22356;
  assign n23688 = ~n23686 & ~n23687;
  assign n23689 = ~n23685 & n23688;
  assign n23690 = n6397 & ~n22556;
  assign n23691 = n23689 & ~n23690;
  assign n23692 =  a[14]  & ~n23691;
  assign n23693 = ~n23691 & ~n23692;
  assign n23694 =  a[14]  & ~n23692;
  assign n23695 = ~n23693 & ~n23694;
  assign n23696 = ~n23619 & ~n23623;
  assign n23697 = ~n23622 & ~n23623;
  assign n23698 = ~n23696 & ~n23697;
  assign n23699 = ~n23695 & ~n23698;
  assign n23700 = ~n23695 & ~n23699;
  assign n23701 = ~n23698 & ~n23699;
  assign n23702 = ~n23700 & ~n23701;
  assign n23703 = n23405 & n23617;
  assign n23704 = ~n23618 & ~n23703;
  assign n23705 = n7101 & n22356;
  assign n23706 = n6402 & n22362;
  assign n23707 = n6951 & n22359;
  assign n23708 = ~n23706 & ~n23707;
  assign n23709 = ~n23705 & n23708;
  assign n23710 = ~n6397 & n23709;
  assign n23711 = n23345 & n23709;
  assign n23712 = ~n23710 & ~n23711;
  assign n23713 =  a[14]  & ~n23712;
  assign n23714 = ~ a[14]  & n23712;
  assign n23715 = ~n23713 & ~n23714;
  assign n23716 = n23704 & ~n23715;
  assign n23717 = n23423 & n23615;
  assign n23718 = ~n23616 & ~n23717;
  assign n23719 = n7101 & n22359;
  assign n23720 = n6402 & n22365;
  assign n23721 = n6951 & n22362;
  assign n23722 = ~n23720 & ~n23721;
  assign n23723 = ~n23719 & n23722;
  assign n23724 = ~n6397 & n23723;
  assign n23725 = ~n23368 & n23723;
  assign n23726 = ~n23724 & ~n23725;
  assign n23727 =  a[14]  & ~n23726;
  assign n23728 = ~ a[14]  & n23726;
  assign n23729 = ~n23727 & ~n23728;
  assign n23730 = n23718 & ~n23729;
  assign n23731 = n23441 & n23613;
  assign n23732 = ~n23614 & ~n23731;
  assign n23733 = n7101 & n22362;
  assign n23734 = n6402 & n22368;
  assign n23735 = n6951 & n22365;
  assign n23736 = ~n23734 & ~n23735;
  assign n23737 = ~n23733 & n23736;
  assign n23738 = ~n6397 & n23737;
  assign n23739 = n23320 & n23737;
  assign n23740 = ~n23738 & ~n23739;
  assign n23741 =  a[14]  & ~n23740;
  assign n23742 = ~ a[14]  & n23740;
  assign n23743 = ~n23741 & ~n23742;
  assign n23744 = n23732 & ~n23743;
  assign n23745 = n7101 & n22365;
  assign n23746 = n6402 & n22371;
  assign n23747 = n6951 & n22368;
  assign n23748 = ~n23746 & ~n23747;
  assign n23749 = ~n23745 & n23748;
  assign n23750 = n6397 & ~n22993;
  assign n23751 = n23749 & ~n23750;
  assign n23752 =  a[14]  & ~n23751;
  assign n23753 = ~n23751 & ~n23752;
  assign n23754 =  a[14]  & ~n23752;
  assign n23755 = ~n23753 & ~n23754;
  assign n23756 = n23609 & ~n23611;
  assign n23757 = ~n23612 & ~n23756;
  assign n23758 = ~n23755 & n23757;
  assign n23759 = ~n23755 & ~n23758;
  assign n23760 = n23757 & ~n23758;
  assign n23761 = ~n23759 & ~n23760;
  assign n23762 = n7101 & n22368;
  assign n23763 = n6402 & n22374;
  assign n23764 = n6951 & n22371;
  assign n23765 = ~n23763 & ~n23764;
  assign n23766 = ~n23762 & n23765;
  assign n23767 = n6397 & n23006;
  assign n23768 = n23766 & ~n23767;
  assign n23769 =  a[14]  & ~n23768;
  assign n23770 = ~n23768 & ~n23769;
  assign n23771 =  a[14]  & ~n23769;
  assign n23772 = ~n23770 & ~n23771;
  assign n23773 = ~n23604 & ~n23608;
  assign n23774 = ~n23607 & ~n23608;
  assign n23775 = ~n23773 & ~n23774;
  assign n23776 = ~n23772 & ~n23775;
  assign n23777 = ~n23772 & ~n23776;
  assign n23778 = ~n23775 & ~n23776;
  assign n23779 = ~n23777 & ~n23778;
  assign n23780 = n7101 & n22371;
  assign n23781 = n6402 & n22377;
  assign n23782 = n6951 & n22374;
  assign n23783 = ~n23781 & ~n23782;
  assign n23784 = ~n23780 & n23783;
  assign n23785 = n6397 & n23025;
  assign n23786 = n23784 & ~n23785;
  assign n23787 =  a[14]  & ~n23786;
  assign n23788 = ~n23786 & ~n23787;
  assign n23789 =  a[14]  & ~n23787;
  assign n23790 = ~n23788 & ~n23789;
  assign n23791 = ~n23599 & ~n23603;
  assign n23792 = ~n23602 & ~n23603;
  assign n23793 = ~n23791 & ~n23792;
  assign n23794 = ~n23790 & ~n23793;
  assign n23795 = ~n23790 & ~n23794;
  assign n23796 = ~n23793 & ~n23794;
  assign n23797 = ~n23795 & ~n23796;
  assign n23798 = n23500 & n23597;
  assign n23799 = ~n23598 & ~n23798;
  assign n23800 = n7101 & n22374;
  assign n23801 = n6402 & n22380;
  assign n23802 = n6951 & n22377;
  assign n23803 = ~n23801 & ~n23802;
  assign n23804 = ~n23800 & n23803;
  assign n23805 = ~n6397 & n23804;
  assign n23806 = ~n22569 & n23804;
  assign n23807 = ~n23805 & ~n23806;
  assign n23808 =  a[14]  & ~n23807;
  assign n23809 = ~ a[14]  & n23807;
  assign n23810 = ~n23808 & ~n23809;
  assign n23811 = n23799 & ~n23810;
  assign n23812 = n23593 & ~n23595;
  assign n23813 = ~n23596 & ~n23812;
  assign n23814 = n7101 & n22377;
  assign n23815 = n6402 & n22384;
  assign n23816 = n6951 & n22380;
  assign n23817 = ~n23815 & ~n23816;
  assign n23818 = ~n23814 & n23817;
  assign n23819 = ~n6397 & n23818;
  assign n23820 = n22834 & n23818;
  assign n23821 = ~n23819 & ~n23820;
  assign n23822 =  a[14]  & ~n23821;
  assign n23823 = ~ a[14]  & n23821;
  assign n23824 = ~n23822 & ~n23823;
  assign n23825 = n23813 & ~n23824;
  assign n23826 = n23532 & n23591;
  assign n23827 = ~n23592 & ~n23826;
  assign n23828 = n7101 & n22380;
  assign n23829 = n6402 & n22387;
  assign n23830 = n6951 & n22384;
  assign n23831 = ~n23829 & ~n23830;
  assign n23832 = ~n23828 & n23831;
  assign n23833 = ~n6397 & n23832;
  assign n23834 = ~n22850 & n23832;
  assign n23835 = ~n23833 & ~n23834;
  assign n23836 =  a[14]  & ~n23835;
  assign n23837 = ~ a[14]  & n23835;
  assign n23838 = ~n23836 & ~n23837;
  assign n23839 = n23827 & ~n23838;
  assign n23840 = n7101 & n22384;
  assign n23841 = n6402 & n22390;
  assign n23842 = n6951 & n22387;
  assign n23843 = ~n23841 & ~n23842;
  assign n23844 = ~n23840 & n23843;
  assign n23845 = n6397 & n22806;
  assign n23846 = n23844 & ~n23845;
  assign n23847 =  a[14]  & ~n23846;
  assign n23848 = ~n23846 & ~n23847;
  assign n23849 =  a[14]  & ~n23847;
  assign n23850 = ~n23848 & ~n23849;
  assign n23851 = n23587 & ~n23589;
  assign n23852 = ~n23590 & ~n23851;
  assign n23853 = ~n23850 & n23852;
  assign n23854 = ~n23850 & ~n23853;
  assign n23855 = n23852 & ~n23853;
  assign n23856 = ~n23854 & ~n23855;
  assign n23857 = ~n23574 & ~n23586;
  assign n23858 = ~n23585 & ~n23586;
  assign n23859 = ~n23857 & ~n23858;
  assign n23860 = n7101 & n22387;
  assign n23861 = n6402 & n22393;
  assign n23862 = n6951 & n22390;
  assign n23863 = ~n23861 & ~n23862;
  assign n23864 = ~n23860 & n23863;
  assign n23865 = ~n6397 & n23864;
  assign n23866 = ~n22582 & n23864;
  assign n23867 = ~n23865 & ~n23866;
  assign n23868 =  a[14]  & ~n23867;
  assign n23869 = ~ a[14]  & n23867;
  assign n23870 = ~n23868 & ~n23869;
  assign n23871 = ~n23859 & ~n23870;
  assign n23872 = n7101 & n22390;
  assign n23873 = n6402 & n22396;
  assign n23874 = n6951 & n22393;
  assign n23875 = ~n23873 & ~n23874;
  assign n23876 = ~n23872 & n23875;
  assign n23877 = n6397 & n22649;
  assign n23878 = n23876 & ~n23877;
  assign n23879 =  a[14]  & ~n23878;
  assign n23880 = ~n23878 & ~n23879;
  assign n23881 =  a[14]  & ~n23879;
  assign n23882 = ~n23880 & ~n23881;
  assign n23883 = ~n23558 & n23569;
  assign n23884 = ~n23570 & ~n23883;
  assign n23885 = ~n23882 & n23884;
  assign n23886 = ~n23882 & ~n23885;
  assign n23887 = n23884 & ~n23885;
  assign n23888 = ~n23886 & ~n23887;
  assign n23889 = n23555 & ~n23557;
  assign n23890 = ~n23558 & ~n23889;
  assign n23891 = n7101 & n22393;
  assign n23892 = n6402 & n22399;
  assign n23893 = n6951 & n22396;
  assign n23894 = ~n23892 & ~n23893;
  assign n23895 = ~n23891 & n23894;
  assign n23896 = ~n6397 & n23895;
  assign n23897 = ~n22671 & n23895;
  assign n23898 = ~n23896 & ~n23897;
  assign n23899 =  a[14]  & ~n23898;
  assign n23900 = ~ a[14]  & n23898;
  assign n23901 = ~n23899 & ~n23900;
  assign n23902 = n23890 & ~n23901;
  assign n23903 = n6951 & ~n22406;
  assign n23904 = n7101 & n22402;
  assign n23905 = ~n23903 & ~n23904;
  assign n23906 = n6397 & ~n22609;
  assign n23907 = n23905 & ~n23906;
  assign n23908 =  a[14]  & ~n23907;
  assign n23909 =  a[14]  & ~n23908;
  assign n23910 = ~n23907 & ~n23908;
  assign n23911 = ~n23909 & ~n23910;
  assign n23912 = ~n6393 & ~n22406;
  assign n23913 =  a[14]  & ~n23912;
  assign n23914 = ~n23911 & n23913;
  assign n23915 = n7101 & n22399;
  assign n23916 = n6402 & ~n22406;
  assign n23917 = n6951 & n22402;
  assign n23918 = ~n23916 & ~n23917;
  assign n23919 = ~n23915 & n23918;
  assign n23920 = ~n6397 & n23919;
  assign n23921 = n22625 & n23919;
  assign n23922 = ~n23920 & ~n23921;
  assign n23923 =  a[14]  & ~n23922;
  assign n23924 = ~ a[14]  & n23922;
  assign n23925 = ~n23923 & ~n23924;
  assign n23926 = n23914 & ~n23925;
  assign n23927 = n23556 & n23926;
  assign n23928 = n23926 & ~n23927;
  assign n23929 = n23556 & ~n23927;
  assign n23930 = ~n23928 & ~n23929;
  assign n23931 = n7101 & n22396;
  assign n23932 = n6402 & n22402;
  assign n23933 = n6951 & n22399;
  assign n23934 = ~n23932 & ~n23933;
  assign n23935 = ~n23931 & n23934;
  assign n23936 = n6397 & n22595;
  assign n23937 = n23935 & ~n23936;
  assign n23938 =  a[14]  & ~n23937;
  assign n23939 =  a[14]  & ~n23938;
  assign n23940 = ~n23937 & ~n23938;
  assign n23941 = ~n23939 & ~n23940;
  assign n23942 = ~n23930 & ~n23941;
  assign n23943 = ~n23927 & ~n23942;
  assign n23944 = ~n23890 & n23901;
  assign n23945 = ~n23902 & ~n23944;
  assign n23946 = ~n23943 & n23945;
  assign n23947 = ~n23902 & ~n23946;
  assign n23948 = ~n23888 & ~n23947;
  assign n23949 = ~n23885 & ~n23948;
  assign n23950 = n23859 & n23870;
  assign n23951 = ~n23871 & ~n23950;
  assign n23952 = ~n23949 & n23951;
  assign n23953 = ~n23871 & ~n23952;
  assign n23954 = ~n23856 & ~n23953;
  assign n23955 = ~n23853 & ~n23954;
  assign n23956 = n23827 & ~n23839;
  assign n23957 = ~n23838 & ~n23839;
  assign n23958 = ~n23956 & ~n23957;
  assign n23959 = ~n23955 & ~n23958;
  assign n23960 = ~n23839 & ~n23959;
  assign n23961 = n23813 & ~n23825;
  assign n23962 = ~n23824 & ~n23825;
  assign n23963 = ~n23961 & ~n23962;
  assign n23964 = ~n23960 & ~n23963;
  assign n23965 = ~n23825 & ~n23964;
  assign n23966 = ~n23799 & n23810;
  assign n23967 = ~n23811 & ~n23966;
  assign n23968 = ~n23965 & n23967;
  assign n23969 = ~n23811 & ~n23968;
  assign n23970 = ~n23797 & ~n23969;
  assign n23971 = ~n23794 & ~n23970;
  assign n23972 = ~n23779 & ~n23971;
  assign n23973 = ~n23776 & ~n23972;
  assign n23974 = ~n23761 & ~n23973;
  assign n23975 = ~n23758 & ~n23974;
  assign n23976 = n23732 & ~n23744;
  assign n23977 = ~n23743 & ~n23744;
  assign n23978 = ~n23976 & ~n23977;
  assign n23979 = ~n23975 & ~n23978;
  assign n23980 = ~n23744 & ~n23979;
  assign n23981 = n23718 & ~n23730;
  assign n23982 = ~n23729 & ~n23730;
  assign n23983 = ~n23981 & ~n23982;
  assign n23984 = ~n23980 & ~n23983;
  assign n23985 = ~n23730 & ~n23984;
  assign n23986 = ~n23704 & n23715;
  assign n23987 = ~n23716 & ~n23986;
  assign n23988 = ~n23985 & n23987;
  assign n23989 = ~n23716 & ~n23988;
  assign n23990 = ~n23702 & ~n23989;
  assign n23991 = ~n23699 & ~n23990;
  assign n23992 = ~n23684 & ~n23991;
  assign n23993 = ~n23681 & ~n23992;
  assign n23994 = n23650 & ~n23665;
  assign n23995 = ~n23664 & ~n23665;
  assign n23996 = ~n23994 & ~n23995;
  assign n23997 = ~n23993 & ~n23996;
  assign n23998 = ~n23665 & ~n23997;
  assign n23999 = n23633 & ~n23648;
  assign n24000 = ~n23647 & ~n23648;
  assign n24001 = ~n23999 & ~n24000;
  assign n24002 = ~n23998 & ~n24001;
  assign n24003 = ~n23648 & ~n24002;
  assign n24004 = n6233 & n22350;
  assign n24005 = n5663 & n22356;
  assign n24006 = n5939 & n22353;
  assign n24007 = ~n24005 & ~n24006;
  assign n24008 = ~n24004 & n24007;
  assign n24009 = n5666 & n23672;
  assign n24010 = n24008 & ~n24009;
  assign n24011 =  a[17]  & ~n24010;
  assign n24012 = ~n24010 & ~n24011;
  assign n24013 =  a[17]  & ~n24011;
  assign n24014 = ~n24012 & ~n24013;
  assign n24015 = ~n23326 & ~n23330;
  assign n24016 = n4694 & n22368;
  assign n24017 = n4533 & n22374;
  assign n24018 = n4604 & n22371;
  assign n24019 = ~n24017 & ~n24018;
  assign n24020 = ~n24016 & n24019;
  assign n24021 = n4536 & n23006;
  assign n24022 = n24020 & ~n24021;
  assign n24023 =  a[23]  & ~n24022;
  assign n24024 = ~n24022 & ~n24023;
  assign n24025 =  a[23]  & ~n24023;
  assign n24026 = ~n24024 & ~n24025;
  assign n24027 = ~n23296 & ~n23300;
  assign n24028 = n3457 & n22387;
  assign n24029 = n3542 & n22393;
  assign n24030 = n3606 & n22390;
  assign n24031 = ~n24029 & ~n24030;
  assign n24032 = ~n24028 & n24031;
  assign n24033 = n3368 & n22582;
  assign n24034 = n24032 & ~n24033;
  assign n24035 =  a[29]  & ~n24034;
  assign n24036 = ~n24034 & ~n24035;
  assign n24037 =  a[29]  & ~n24035;
  assign n24038 = ~n24036 & ~n24037;
  assign n24039 = ~n23270 & ~n23273;
  assign n24040 = n116 & ~n511;
  assign n24041 = ~n514 & n24040;
  assign n24042 = n1971 & n5002;
  assign n24043 = n24041 & n24042;
  assign n24044 = n4216 & n24043;
  assign n24045 = n1621 & n24044;
  assign n24046 = n5296 & n24045;
  assign n24047 = n916 & n24046;
  assign n24048 = n3290 & n24047;
  assign n24049 = n2346 & n24048;
  assign n24050 = n291 & n24049;
  assign n24051 = n471 & n24050;
  assign n24052 = n1531 & n24051;
  assign n24053 = n520 & n24052;
  assign n24054 = ~n118 & n24053;
  assign n24055 = ~n102 & n24054;
  assign n24056 = ~n791 & n24055;
  assign n24057 = ~n225 & n24056;
  assign n24058 = n3020 & n22396;
  assign n24059 = n3028 & n22399;
  assign n24060 = n3023 & n22402;
  assign n24061 = n75 & n22595;
  assign n24062 = ~n24060 & ~n24061;
  assign n24063 = ~n24059 & n24062;
  assign n24064 = ~n24058 & n24063;
  assign n24065 = ~n24057 & ~n24064;
  assign n24066 = ~n24057 & ~n24065;
  assign n24067 = ~n24064 & ~n24065;
  assign n24068 = ~n24066 & ~n24067;
  assign n24069 = ~n24039 & ~n24068;
  assign n24070 = ~n24039 & ~n24069;
  assign n24071 = ~n24068 & ~n24069;
  assign n24072 = ~n24070 & ~n24071;
  assign n24073 = ~n24038 & ~n24072;
  assign n24074 = ~n24038 & ~n24073;
  assign n24075 = ~n24072 & ~n24073;
  assign n24076 = ~n24074 & ~n24075;
  assign n24077 = ~n23277 & ~n23283;
  assign n24078 = n24076 & n24077;
  assign n24079 = ~n24076 & ~n24077;
  assign n24080 = ~n24078 & ~n24079;
  assign n24081 = n3884 & n22377;
  assign n24082 = n3967 & n22384;
  assign n24083 = n4046 & n22380;
  assign n24084 = ~n24082 & ~n24083;
  assign n24085 = ~n24081 & n24084;
  assign n24086 = ~n4050 & n24085;
  assign n24087 = n22834 & n24085;
  assign n24088 = ~n24086 & ~n24087;
  assign n24089 =  a[26]  & ~n24088;
  assign n24090 = ~ a[26]  & n24088;
  assign n24091 = ~n24089 & ~n24090;
  assign n24092 = n24080 & ~n24091;
  assign n24093 = n24080 & ~n24092;
  assign n24094 = ~n24091 & ~n24092;
  assign n24095 = ~n24093 & ~n24094;
  assign n24096 = ~n24027 & ~n24095;
  assign n24097 = ~n24027 & ~n24096;
  assign n24098 = ~n24095 & ~n24096;
  assign n24099 = ~n24097 & ~n24098;
  assign n24100 = ~n24026 & ~n24099;
  assign n24101 = ~n24026 & ~n24100;
  assign n24102 = ~n24099 & ~n24100;
  assign n24103 = ~n24101 & ~n24102;
  assign n24104 = ~n23304 & ~n23310;
  assign n24105 = n24103 & n24104;
  assign n24106 = ~n24103 & ~n24104;
  assign n24107 = ~n24105 & ~n24106;
  assign n24108 = n5496 & n22359;
  assign n24109 = n4935 & n22365;
  assign n24110 = n5407 & n22362;
  assign n24111 = ~n24109 & ~n24110;
  assign n24112 = ~n24108 & n24111;
  assign n24113 = ~n4938 & n24112;
  assign n24114 = ~n23368 & n24112;
  assign n24115 = ~n24113 & ~n24114;
  assign n24116 =  a[20]  & ~n24115;
  assign n24117 = ~ a[20]  & n24115;
  assign n24118 = ~n24116 & ~n24117;
  assign n24119 = n24107 & ~n24118;
  assign n24120 = n24107 & ~n24119;
  assign n24121 = ~n24118 & ~n24119;
  assign n24122 = ~n24120 & ~n24121;
  assign n24123 = ~n24015 & ~n24122;
  assign n24124 = ~n24015 & ~n24123;
  assign n24125 = ~n24122 & ~n24123;
  assign n24126 = ~n24124 & ~n24125;
  assign n24127 = ~n24014 & ~n24126;
  assign n24128 = ~n24014 & ~n24127;
  assign n24129 = ~n24126 & ~n24127;
  assign n24130 = ~n24128 & ~n24129;
  assign n24131 = ~n23334 & ~n23632;
  assign n24132 = n24130 & n24131;
  assign n24133 = ~n24130 & ~n24131;
  assign n24134 = ~n24132 & ~n24133;
  assign n24135 = n7101 & n22341;
  assign n24136 = n6402 & n22347;
  assign n24137 = n6951 & n22344;
  assign n24138 = ~n24136 & ~n24137;
  assign n24139 = ~n24135 & n24138;
  assign n24140 = ~n6397 & n24139;
  assign n24141 = n22480 & ~n22482;
  assign n24142 = ~n22483 & ~n24141;
  assign n24143 = n24139 & ~n24142;
  assign n24144 = ~n24140 & ~n24143;
  assign n24145 =  a[14]  & ~n24144;
  assign n24146 = ~ a[14]  & n24144;
  assign n24147 = ~n24145 & ~n24146;
  assign n24148 = n24134 & ~n24147;
  assign n24149 = n24134 & ~n24148;
  assign n24150 = ~n24147 & ~n24148;
  assign n24151 = ~n24149 & ~n24150;
  assign n24152 = ~n24003 & ~n24151;
  assign n24153 = ~n24003 & ~n24152;
  assign n24154 = ~n24151 & ~n24152;
  assign n24155 = ~n24153 & ~n24154;
  assign n24156 = ~n22548 & ~n24155;
  assign n24157 = ~n22548 & ~n24156;
  assign n24158 = ~n24155 & ~n24156;
  assign n24159 = ~n24157 & ~n24158;
  assign n24160 = n7983 & n22335;
  assign n24161 = n7291 & n22341;
  assign n24162 = n7632 & n22338;
  assign n24163 = ~n24161 & ~n24162;
  assign n24164 = ~n24160 & n24163;
  assign n24165 = ~n22488 & ~n22491;
  assign n24166 = ~n22489 & n22492;
  assign n24167 = ~n24165 & ~n24166;
  assign n24168 = n7294 & ~n24167;
  assign n24169 = n24164 & ~n24168;
  assign n24170 =  a[11]  & ~n24169;
  assign n24171 = ~n24169 & ~n24170;
  assign n24172 =  a[11]  & ~n24170;
  assign n24173 = ~n24171 & ~n24172;
  assign n24174 = ~n23998 & ~n24002;
  assign n24175 = ~n24001 & ~n24002;
  assign n24176 = ~n24174 & ~n24175;
  assign n24177 = ~n24173 & ~n24176;
  assign n24178 = ~n24173 & ~n24177;
  assign n24179 = ~n24176 & ~n24177;
  assign n24180 = ~n24178 & ~n24179;
  assign n24181 = n7983 & n22338;
  assign n24182 = n7291 & n22344;
  assign n24183 = n7632 & n22341;
  assign n24184 = ~n24182 & ~n24183;
  assign n24185 = ~n24181 & n24184;
  assign n24186 = ~n22484 & ~n22487;
  assign n24187 = ~n22485 & n22488;
  assign n24188 = ~n24186 & ~n24187;
  assign n24189 = n7294 & ~n24188;
  assign n24190 = n24185 & ~n24189;
  assign n24191 =  a[11]  & ~n24190;
  assign n24192 = ~n24190 & ~n24191;
  assign n24193 =  a[11]  & ~n24191;
  assign n24194 = ~n24192 & ~n24193;
  assign n24195 = ~n23993 & ~n23997;
  assign n24196 = ~n23996 & ~n23997;
  assign n24197 = ~n24195 & ~n24196;
  assign n24198 = ~n24194 & ~n24197;
  assign n24199 = ~n24194 & ~n24198;
  assign n24200 = ~n24197 & ~n24198;
  assign n24201 = ~n24199 & ~n24200;
  assign n24202 = n23684 & n23991;
  assign n24203 = ~n23992 & ~n24202;
  assign n24204 = n7983 & n22341;
  assign n24205 = n7291 & n22347;
  assign n24206 = n7632 & n22344;
  assign n24207 = ~n24205 & ~n24206;
  assign n24208 = ~n24204 & n24207;
  assign n24209 = ~n7294 & n24208;
  assign n24210 = ~n24142 & n24208;
  assign n24211 = ~n24209 & ~n24210;
  assign n24212 =  a[11]  & ~n24211;
  assign n24213 = ~ a[11]  & n24211;
  assign n24214 = ~n24212 & ~n24213;
  assign n24215 = n24203 & ~n24214;
  assign n24216 = n23702 & n23989;
  assign n24217 = ~n23990 & ~n24216;
  assign n24218 = n7983 & n22344;
  assign n24219 = n7291 & n22350;
  assign n24220 = n7632 & n22347;
  assign n24221 = ~n24219 & ~n24220;
  assign n24222 = ~n24218 & n24221;
  assign n24223 = ~n7294 & n24222;
  assign n24224 = n23642 & n24222;
  assign n24225 = ~n24223 & ~n24224;
  assign n24226 =  a[11]  & ~n24225;
  assign n24227 = ~ a[11]  & n24225;
  assign n24228 = ~n24226 & ~n24227;
  assign n24229 = n24217 & ~n24228;
  assign n24230 = n7983 & n22347;
  assign n24231 = n7291 & n22353;
  assign n24232 = n7632 & n22350;
  assign n24233 = ~n24231 & ~n24232;
  assign n24234 = ~n24230 & n24233;
  assign n24235 = n7294 & ~n23659;
  assign n24236 = n24234 & ~n24235;
  assign n24237 =  a[11]  & ~n24236;
  assign n24238 = ~n24236 & ~n24237;
  assign n24239 =  a[11]  & ~n24237;
  assign n24240 = ~n24238 & ~n24239;
  assign n24241 = n23985 & ~n23987;
  assign n24242 = ~n23988 & ~n24241;
  assign n24243 = ~n24240 & n24242;
  assign n24244 = ~n24240 & ~n24243;
  assign n24245 = n24242 & ~n24243;
  assign n24246 = ~n24244 & ~n24245;
  assign n24247 = n7983 & n22350;
  assign n24248 = n7291 & n22356;
  assign n24249 = n7632 & n22353;
  assign n24250 = ~n24248 & ~n24249;
  assign n24251 = ~n24247 & n24250;
  assign n24252 = n7294 & n23672;
  assign n24253 = n24251 & ~n24252;
  assign n24254 =  a[11]  & ~n24253;
  assign n24255 = ~n24253 & ~n24254;
  assign n24256 =  a[11]  & ~n24254;
  assign n24257 = ~n24255 & ~n24256;
  assign n24258 = ~n23980 & ~n23984;
  assign n24259 = ~n23983 & ~n23984;
  assign n24260 = ~n24258 & ~n24259;
  assign n24261 = ~n24257 & ~n24260;
  assign n24262 = ~n24257 & ~n24261;
  assign n24263 = ~n24260 & ~n24261;
  assign n24264 = ~n24262 & ~n24263;
  assign n24265 = n7983 & n22353;
  assign n24266 = n7291 & n22359;
  assign n24267 = n7632 & n22356;
  assign n24268 = ~n24266 & ~n24267;
  assign n24269 = ~n24265 & n24268;
  assign n24270 = n7294 & ~n22556;
  assign n24271 = n24269 & ~n24270;
  assign n24272 =  a[11]  & ~n24271;
  assign n24273 = ~n24271 & ~n24272;
  assign n24274 =  a[11]  & ~n24272;
  assign n24275 = ~n24273 & ~n24274;
  assign n24276 = ~n23975 & ~n23979;
  assign n24277 = ~n23978 & ~n23979;
  assign n24278 = ~n24276 & ~n24277;
  assign n24279 = ~n24275 & ~n24278;
  assign n24280 = ~n24275 & ~n24279;
  assign n24281 = ~n24278 & ~n24279;
  assign n24282 = ~n24280 & ~n24281;
  assign n24283 = n23761 & n23973;
  assign n24284 = ~n23974 & ~n24283;
  assign n24285 = n7983 & n22356;
  assign n24286 = n7291 & n22362;
  assign n24287 = n7632 & n22359;
  assign n24288 = ~n24286 & ~n24287;
  assign n24289 = ~n24285 & n24288;
  assign n24290 = ~n7294 & n24289;
  assign n24291 = n23345 & n24289;
  assign n24292 = ~n24290 & ~n24291;
  assign n24293 =  a[11]  & ~n24292;
  assign n24294 = ~ a[11]  & n24292;
  assign n24295 = ~n24293 & ~n24294;
  assign n24296 = n24284 & ~n24295;
  assign n24297 = n23779 & n23971;
  assign n24298 = ~n23972 & ~n24297;
  assign n24299 = n7983 & n22359;
  assign n24300 = n7291 & n22365;
  assign n24301 = n7632 & n22362;
  assign n24302 = ~n24300 & ~n24301;
  assign n24303 = ~n24299 & n24302;
  assign n24304 = ~n7294 & n24303;
  assign n24305 = ~n23368 & n24303;
  assign n24306 = ~n24304 & ~n24305;
  assign n24307 =  a[11]  & ~n24306;
  assign n24308 = ~ a[11]  & n24306;
  assign n24309 = ~n24307 & ~n24308;
  assign n24310 = n24298 & ~n24309;
  assign n24311 = n23797 & n23969;
  assign n24312 = ~n23970 & ~n24311;
  assign n24313 = n7983 & n22362;
  assign n24314 = n7291 & n22368;
  assign n24315 = n7632 & n22365;
  assign n24316 = ~n24314 & ~n24315;
  assign n24317 = ~n24313 & n24316;
  assign n24318 = ~n7294 & n24317;
  assign n24319 = n23320 & n24317;
  assign n24320 = ~n24318 & ~n24319;
  assign n24321 =  a[11]  & ~n24320;
  assign n24322 = ~ a[11]  & n24320;
  assign n24323 = ~n24321 & ~n24322;
  assign n24324 = n24312 & ~n24323;
  assign n24325 = n7983 & n22365;
  assign n24326 = n7291 & n22371;
  assign n24327 = n7632 & n22368;
  assign n24328 = ~n24326 & ~n24327;
  assign n24329 = ~n24325 & n24328;
  assign n24330 = n7294 & ~n22993;
  assign n24331 = n24329 & ~n24330;
  assign n24332 =  a[11]  & ~n24331;
  assign n24333 = ~n24331 & ~n24332;
  assign n24334 =  a[11]  & ~n24332;
  assign n24335 = ~n24333 & ~n24334;
  assign n24336 = n23965 & ~n23967;
  assign n24337 = ~n23968 & ~n24336;
  assign n24338 = ~n24335 & n24337;
  assign n24339 = ~n24335 & ~n24338;
  assign n24340 = n24337 & ~n24338;
  assign n24341 = ~n24339 & ~n24340;
  assign n24342 = n7983 & n22368;
  assign n24343 = n7291 & n22374;
  assign n24344 = n7632 & n22371;
  assign n24345 = ~n24343 & ~n24344;
  assign n24346 = ~n24342 & n24345;
  assign n24347 = n7294 & n23006;
  assign n24348 = n24346 & ~n24347;
  assign n24349 =  a[11]  & ~n24348;
  assign n24350 = ~n24348 & ~n24349;
  assign n24351 =  a[11]  & ~n24349;
  assign n24352 = ~n24350 & ~n24351;
  assign n24353 = ~n23960 & ~n23964;
  assign n24354 = ~n23963 & ~n23964;
  assign n24355 = ~n24353 & ~n24354;
  assign n24356 = ~n24352 & ~n24355;
  assign n24357 = ~n24352 & ~n24356;
  assign n24358 = ~n24355 & ~n24356;
  assign n24359 = ~n24357 & ~n24358;
  assign n24360 = n7983 & n22371;
  assign n24361 = n7291 & n22377;
  assign n24362 = n7632 & n22374;
  assign n24363 = ~n24361 & ~n24362;
  assign n24364 = ~n24360 & n24363;
  assign n24365 = n7294 & n23025;
  assign n24366 = n24364 & ~n24365;
  assign n24367 =  a[11]  & ~n24366;
  assign n24368 = ~n24366 & ~n24367;
  assign n24369 =  a[11]  & ~n24367;
  assign n24370 = ~n24368 & ~n24369;
  assign n24371 = ~n23955 & ~n23959;
  assign n24372 = ~n23958 & ~n23959;
  assign n24373 = ~n24371 & ~n24372;
  assign n24374 = ~n24370 & ~n24373;
  assign n24375 = ~n24370 & ~n24374;
  assign n24376 = ~n24373 & ~n24374;
  assign n24377 = ~n24375 & ~n24376;
  assign n24378 = n23856 & n23953;
  assign n24379 = ~n23954 & ~n24378;
  assign n24380 = n7983 & n22374;
  assign n24381 = n7291 & n22380;
  assign n24382 = n7632 & n22377;
  assign n24383 = ~n24381 & ~n24382;
  assign n24384 = ~n24380 & n24383;
  assign n24385 = ~n7294 & n24384;
  assign n24386 = ~n22569 & n24384;
  assign n24387 = ~n24385 & ~n24386;
  assign n24388 =  a[11]  & ~n24387;
  assign n24389 = ~ a[11]  & n24387;
  assign n24390 = ~n24388 & ~n24389;
  assign n24391 = n24379 & ~n24390;
  assign n24392 = n23949 & ~n23951;
  assign n24393 = ~n23952 & ~n24392;
  assign n24394 = n7983 & n22377;
  assign n24395 = n7291 & n22384;
  assign n24396 = n7632 & n22380;
  assign n24397 = ~n24395 & ~n24396;
  assign n24398 = ~n24394 & n24397;
  assign n24399 = ~n7294 & n24398;
  assign n24400 = n22834 & n24398;
  assign n24401 = ~n24399 & ~n24400;
  assign n24402 =  a[11]  & ~n24401;
  assign n24403 = ~ a[11]  & n24401;
  assign n24404 = ~n24402 & ~n24403;
  assign n24405 = n24393 & ~n24404;
  assign n24406 = n23888 & n23947;
  assign n24407 = ~n23948 & ~n24406;
  assign n24408 = n7983 & n22380;
  assign n24409 = n7291 & n22387;
  assign n24410 = n7632 & n22384;
  assign n24411 = ~n24409 & ~n24410;
  assign n24412 = ~n24408 & n24411;
  assign n24413 = ~n7294 & n24412;
  assign n24414 = ~n22850 & n24412;
  assign n24415 = ~n24413 & ~n24414;
  assign n24416 =  a[11]  & ~n24415;
  assign n24417 = ~ a[11]  & n24415;
  assign n24418 = ~n24416 & ~n24417;
  assign n24419 = n24407 & ~n24418;
  assign n24420 = n7983 & n22384;
  assign n24421 = n7291 & n22390;
  assign n24422 = n7632 & n22387;
  assign n24423 = ~n24421 & ~n24422;
  assign n24424 = ~n24420 & n24423;
  assign n24425 = n7294 & n22806;
  assign n24426 = n24424 & ~n24425;
  assign n24427 =  a[11]  & ~n24426;
  assign n24428 = ~n24426 & ~n24427;
  assign n24429 =  a[11]  & ~n24427;
  assign n24430 = ~n24428 & ~n24429;
  assign n24431 = n23943 & ~n23945;
  assign n24432 = ~n23946 & ~n24431;
  assign n24433 = ~n24430 & n24432;
  assign n24434 = ~n24430 & ~n24433;
  assign n24435 = n24432 & ~n24433;
  assign n24436 = ~n24434 & ~n24435;
  assign n24437 = ~n23930 & ~n23942;
  assign n24438 = ~n23941 & ~n23942;
  assign n24439 = ~n24437 & ~n24438;
  assign n24440 = n7983 & n22387;
  assign n24441 = n7291 & n22393;
  assign n24442 = n7632 & n22390;
  assign n24443 = ~n24441 & ~n24442;
  assign n24444 = ~n24440 & n24443;
  assign n24445 = ~n7294 & n24444;
  assign n24446 = ~n22582 & n24444;
  assign n24447 = ~n24445 & ~n24446;
  assign n24448 =  a[11]  & ~n24447;
  assign n24449 = ~ a[11]  & n24447;
  assign n24450 = ~n24448 & ~n24449;
  assign n24451 = ~n24439 & ~n24450;
  assign n24452 = n7983 & n22390;
  assign n24453 = n7291 & n22396;
  assign n24454 = n7632 & n22393;
  assign n24455 = ~n24453 & ~n24454;
  assign n24456 = ~n24452 & n24455;
  assign n24457 = n7294 & n22649;
  assign n24458 = n24456 & ~n24457;
  assign n24459 =  a[11]  & ~n24458;
  assign n24460 = ~n24458 & ~n24459;
  assign n24461 =  a[11]  & ~n24459;
  assign n24462 = ~n24460 & ~n24461;
  assign n24463 = ~n23914 & n23925;
  assign n24464 = ~n23926 & ~n24463;
  assign n24465 = ~n24462 & n24464;
  assign n24466 = ~n24462 & ~n24465;
  assign n24467 = n24464 & ~n24465;
  assign n24468 = ~n24466 & ~n24467;
  assign n24469 = n23911 & ~n23913;
  assign n24470 = ~n23914 & ~n24469;
  assign n24471 = n7983 & n22393;
  assign n24472 = n7291 & n22399;
  assign n24473 = n7632 & n22396;
  assign n24474 = ~n24472 & ~n24473;
  assign n24475 = ~n24471 & n24474;
  assign n24476 = ~n7294 & n24475;
  assign n24477 = ~n22671 & n24475;
  assign n24478 = ~n24476 & ~n24477;
  assign n24479 =  a[11]  & ~n24478;
  assign n24480 = ~ a[11]  & n24478;
  assign n24481 = ~n24479 & ~n24480;
  assign n24482 = n24470 & ~n24481;
  assign n24483 = n7632 & ~n22406;
  assign n24484 = n7983 & n22402;
  assign n24485 = ~n24483 & ~n24484;
  assign n24486 = n7294 & ~n22609;
  assign n24487 = n24485 & ~n24486;
  assign n24488 =  a[11]  & ~n24487;
  assign n24489 =  a[11]  & ~n24488;
  assign n24490 = ~n24487 & ~n24488;
  assign n24491 = ~n24489 & ~n24490;
  assign n24492 = ~n7289 & ~n22406;
  assign n24493 =  a[11]  & ~n24492;
  assign n24494 = ~n24491 & n24493;
  assign n24495 = n7983 & n22399;
  assign n24496 = n7291 & ~n22406;
  assign n24497 = n7632 & n22402;
  assign n24498 = ~n24496 & ~n24497;
  assign n24499 = ~n24495 & n24498;
  assign n24500 = ~n7294 & n24499;
  assign n24501 = n22625 & n24499;
  assign n24502 = ~n24500 & ~n24501;
  assign n24503 =  a[11]  & ~n24502;
  assign n24504 = ~ a[11]  & n24502;
  assign n24505 = ~n24503 & ~n24504;
  assign n24506 = n24494 & ~n24505;
  assign n24507 = n23912 & n24506;
  assign n24508 = n24506 & ~n24507;
  assign n24509 = n23912 & ~n24507;
  assign n24510 = ~n24508 & ~n24509;
  assign n24511 = n7983 & n22396;
  assign n24512 = n7291 & n22402;
  assign n24513 = n7632 & n22399;
  assign n24514 = ~n24512 & ~n24513;
  assign n24515 = ~n24511 & n24514;
  assign n24516 = n7294 & n22595;
  assign n24517 = n24515 & ~n24516;
  assign n24518 =  a[11]  & ~n24517;
  assign n24519 =  a[11]  & ~n24518;
  assign n24520 = ~n24517 & ~n24518;
  assign n24521 = ~n24519 & ~n24520;
  assign n24522 = ~n24510 & ~n24521;
  assign n24523 = ~n24507 & ~n24522;
  assign n24524 = ~n24470 & n24481;
  assign n24525 = ~n24482 & ~n24524;
  assign n24526 = ~n24523 & n24525;
  assign n24527 = ~n24482 & ~n24526;
  assign n24528 = ~n24468 & ~n24527;
  assign n24529 = ~n24465 & ~n24528;
  assign n24530 = n24439 & n24450;
  assign n24531 = ~n24451 & ~n24530;
  assign n24532 = ~n24529 & n24531;
  assign n24533 = ~n24451 & ~n24532;
  assign n24534 = ~n24436 & ~n24533;
  assign n24535 = ~n24433 & ~n24534;
  assign n24536 = n24407 & ~n24419;
  assign n24537 = ~n24418 & ~n24419;
  assign n24538 = ~n24536 & ~n24537;
  assign n24539 = ~n24535 & ~n24538;
  assign n24540 = ~n24419 & ~n24539;
  assign n24541 = n24393 & ~n24405;
  assign n24542 = ~n24404 & ~n24405;
  assign n24543 = ~n24541 & ~n24542;
  assign n24544 = ~n24540 & ~n24543;
  assign n24545 = ~n24405 & ~n24544;
  assign n24546 = ~n24379 & n24390;
  assign n24547 = ~n24391 & ~n24546;
  assign n24548 = ~n24545 & n24547;
  assign n24549 = ~n24391 & ~n24548;
  assign n24550 = ~n24377 & ~n24549;
  assign n24551 = ~n24374 & ~n24550;
  assign n24552 = ~n24359 & ~n24551;
  assign n24553 = ~n24356 & ~n24552;
  assign n24554 = ~n24341 & ~n24553;
  assign n24555 = ~n24338 & ~n24554;
  assign n24556 = n24312 & ~n24324;
  assign n24557 = ~n24323 & ~n24324;
  assign n24558 = ~n24556 & ~n24557;
  assign n24559 = ~n24555 & ~n24558;
  assign n24560 = ~n24324 & ~n24559;
  assign n24561 = n24298 & ~n24310;
  assign n24562 = ~n24309 & ~n24310;
  assign n24563 = ~n24561 & ~n24562;
  assign n24564 = ~n24560 & ~n24563;
  assign n24565 = ~n24310 & ~n24564;
  assign n24566 = ~n24284 & n24295;
  assign n24567 = ~n24296 & ~n24566;
  assign n24568 = ~n24565 & n24567;
  assign n24569 = ~n24296 & ~n24568;
  assign n24570 = ~n24282 & ~n24569;
  assign n24571 = ~n24279 & ~n24570;
  assign n24572 = ~n24264 & ~n24571;
  assign n24573 = ~n24261 & ~n24572;
  assign n24574 = ~n24246 & ~n24573;
  assign n24575 = ~n24243 & ~n24574;
  assign n24576 = n24217 & ~n24229;
  assign n24577 = ~n24228 & ~n24229;
  assign n24578 = ~n24576 & ~n24577;
  assign n24579 = ~n24575 & ~n24578;
  assign n24580 = ~n24229 & ~n24579;
  assign n24581 = ~n24203 & n24214;
  assign n24582 = ~n24215 & ~n24581;
  assign n24583 = ~n24580 & n24582;
  assign n24584 = ~n24215 & ~n24583;
  assign n24585 = ~n24201 & ~n24584;
  assign n24586 = ~n24198 & ~n24585;
  assign n24587 = ~n24180 & ~n24586;
  assign n24588 = ~n24177 & ~n24587;
  assign n24589 = n24159 & n24588;
  assign n24590 = ~n24159 & ~n24588;
  assign n24591 = ~n24589 & ~n24590;
  assign n24592 = n9331 & n22323;
  assign n24593 = n8418 & n22329;
  assign n24594 = n8860 & n22326;
  assign n24595 = ~n24593 & ~n24594;
  assign n24596 = ~n24592 & n24595;
  assign n24597 = ~n8421 & n24596;
  assign n24598 = n22504 & ~n22506;
  assign n24599 = ~n22507 & ~n24598;
  assign n24600 = n24596 & ~n24599;
  assign n24601 = ~n24597 & ~n24600;
  assign n24602 =  a[8]  & ~n24601;
  assign n24603 = ~ a[8]  & n24601;
  assign n24604 = ~n24602 & ~n24603;
  assign n24605 = n24591 & ~n24604;
  assign n24606 = n24180 & n24586;
  assign n24607 = ~n24587 & ~n24606;
  assign n24608 = n9331 & n22326;
  assign n24609 = n8418 & n22332;
  assign n24610 = n8860 & n22329;
  assign n24611 = ~n24609 & ~n24610;
  assign n24612 = ~n24608 & n24611;
  assign n24613 = ~n8421 & n24612;
  assign n24614 = ~n22500 & ~n22503;
  assign n24615 = ~n22501 & n22504;
  assign n24616 = ~n24614 & ~n24615;
  assign n24617 = n24612 & n24616;
  assign n24618 = ~n24613 & ~n24617;
  assign n24619 =  a[8]  & ~n24618;
  assign n24620 = ~ a[8]  & n24618;
  assign n24621 = ~n24619 & ~n24620;
  assign n24622 = n24607 & ~n24621;
  assign n24623 = n24201 & n24584;
  assign n24624 = ~n24585 & ~n24623;
  assign n24625 = n9331 & n22329;
  assign n24626 = n8418 & n22335;
  assign n24627 = n8860 & n22332;
  assign n24628 = ~n24626 & ~n24627;
  assign n24629 = ~n24625 & n24628;
  assign n24630 = ~n8421 & n24629;
  assign n24631 = ~n22496 & ~n22499;
  assign n24632 = ~n22497 & n22500;
  assign n24633 = ~n24631 & ~n24632;
  assign n24634 = n24629 & n24633;
  assign n24635 = ~n24630 & ~n24634;
  assign n24636 =  a[8]  & ~n24635;
  assign n24637 = ~ a[8]  & n24635;
  assign n24638 = ~n24636 & ~n24637;
  assign n24639 = n24624 & ~n24638;
  assign n24640 = n9331 & n22332;
  assign n24641 = n8418 & n22338;
  assign n24642 = n8860 & n22335;
  assign n24643 = ~n24641 & ~n24642;
  assign n24644 = ~n24640 & n24643;
  assign n24645 = n8421 & n22542;
  assign n24646 = n24644 & ~n24645;
  assign n24647 =  a[8]  & ~n24646;
  assign n24648 = ~n24646 & ~n24647;
  assign n24649 =  a[8]  & ~n24647;
  assign n24650 = ~n24648 & ~n24649;
  assign n24651 = n24580 & ~n24582;
  assign n24652 = ~n24583 & ~n24651;
  assign n24653 = ~n24650 & n24652;
  assign n24654 = ~n24650 & ~n24653;
  assign n24655 = n24652 & ~n24653;
  assign n24656 = ~n24654 & ~n24655;
  assign n24657 = n9331 & n22335;
  assign n24658 = n8418 & n22341;
  assign n24659 = n8860 & n22338;
  assign n24660 = ~n24658 & ~n24659;
  assign n24661 = ~n24657 & n24660;
  assign n24662 = n8421 & ~n24167;
  assign n24663 = n24661 & ~n24662;
  assign n24664 =  a[8]  & ~n24663;
  assign n24665 = ~n24663 & ~n24664;
  assign n24666 =  a[8]  & ~n24664;
  assign n24667 = ~n24665 & ~n24666;
  assign n24668 = ~n24575 & ~n24579;
  assign n24669 = ~n24578 & ~n24579;
  assign n24670 = ~n24668 & ~n24669;
  assign n24671 = ~n24667 & ~n24670;
  assign n24672 = ~n24667 & ~n24671;
  assign n24673 = ~n24670 & ~n24671;
  assign n24674 = ~n24672 & ~n24673;
  assign n24675 = n24246 & n24573;
  assign n24676 = ~n24574 & ~n24675;
  assign n24677 = n9331 & n22338;
  assign n24678 = n8418 & n22344;
  assign n24679 = n8860 & n22341;
  assign n24680 = ~n24678 & ~n24679;
  assign n24681 = ~n24677 & n24680;
  assign n24682 = ~n8421 & n24681;
  assign n24683 = n24188 & n24681;
  assign n24684 = ~n24682 & ~n24683;
  assign n24685 =  a[8]  & ~n24684;
  assign n24686 = ~ a[8]  & n24684;
  assign n24687 = ~n24685 & ~n24686;
  assign n24688 = n24676 & ~n24687;
  assign n24689 = n24264 & n24571;
  assign n24690 = ~n24572 & ~n24689;
  assign n24691 = n9331 & n22341;
  assign n24692 = n8418 & n22347;
  assign n24693 = n8860 & n22344;
  assign n24694 = ~n24692 & ~n24693;
  assign n24695 = ~n24691 & n24694;
  assign n24696 = ~n8421 & n24695;
  assign n24697 = ~n24142 & n24695;
  assign n24698 = ~n24696 & ~n24697;
  assign n24699 =  a[8]  & ~n24698;
  assign n24700 = ~ a[8]  & n24698;
  assign n24701 = ~n24699 & ~n24700;
  assign n24702 = n24690 & ~n24701;
  assign n24703 = n24282 & n24569;
  assign n24704 = ~n24570 & ~n24703;
  assign n24705 = n9331 & n22344;
  assign n24706 = n8418 & n22350;
  assign n24707 = n8860 & n22347;
  assign n24708 = ~n24706 & ~n24707;
  assign n24709 = ~n24705 & n24708;
  assign n24710 = ~n8421 & n24709;
  assign n24711 = n23642 & n24709;
  assign n24712 = ~n24710 & ~n24711;
  assign n24713 =  a[8]  & ~n24712;
  assign n24714 = ~ a[8]  & n24712;
  assign n24715 = ~n24713 & ~n24714;
  assign n24716 = n24704 & ~n24715;
  assign n24717 = n9331 & n22347;
  assign n24718 = n8418 & n22353;
  assign n24719 = n8860 & n22350;
  assign n24720 = ~n24718 & ~n24719;
  assign n24721 = ~n24717 & n24720;
  assign n24722 = n8421 & ~n23659;
  assign n24723 = n24721 & ~n24722;
  assign n24724 =  a[8]  & ~n24723;
  assign n24725 = ~n24723 & ~n24724;
  assign n24726 =  a[8]  & ~n24724;
  assign n24727 = ~n24725 & ~n24726;
  assign n24728 = n24565 & ~n24567;
  assign n24729 = ~n24568 & ~n24728;
  assign n24730 = ~n24727 & n24729;
  assign n24731 = ~n24727 & ~n24730;
  assign n24732 = n24729 & ~n24730;
  assign n24733 = ~n24731 & ~n24732;
  assign n24734 = n9331 & n22350;
  assign n24735 = n8418 & n22356;
  assign n24736 = n8860 & n22353;
  assign n24737 = ~n24735 & ~n24736;
  assign n24738 = ~n24734 & n24737;
  assign n24739 = n8421 & n23672;
  assign n24740 = n24738 & ~n24739;
  assign n24741 =  a[8]  & ~n24740;
  assign n24742 = ~n24740 & ~n24741;
  assign n24743 =  a[8]  & ~n24741;
  assign n24744 = ~n24742 & ~n24743;
  assign n24745 = ~n24560 & ~n24564;
  assign n24746 = ~n24563 & ~n24564;
  assign n24747 = ~n24745 & ~n24746;
  assign n24748 = ~n24744 & ~n24747;
  assign n24749 = ~n24744 & ~n24748;
  assign n24750 = ~n24747 & ~n24748;
  assign n24751 = ~n24749 & ~n24750;
  assign n24752 = n9331 & n22353;
  assign n24753 = n8418 & n22359;
  assign n24754 = n8860 & n22356;
  assign n24755 = ~n24753 & ~n24754;
  assign n24756 = ~n24752 & n24755;
  assign n24757 = n8421 & ~n22556;
  assign n24758 = n24756 & ~n24757;
  assign n24759 =  a[8]  & ~n24758;
  assign n24760 = ~n24758 & ~n24759;
  assign n24761 =  a[8]  & ~n24759;
  assign n24762 = ~n24760 & ~n24761;
  assign n24763 = ~n24555 & ~n24559;
  assign n24764 = ~n24558 & ~n24559;
  assign n24765 = ~n24763 & ~n24764;
  assign n24766 = ~n24762 & ~n24765;
  assign n24767 = ~n24762 & ~n24766;
  assign n24768 = ~n24765 & ~n24766;
  assign n24769 = ~n24767 & ~n24768;
  assign n24770 = n24341 & n24553;
  assign n24771 = ~n24554 & ~n24770;
  assign n24772 = n9331 & n22356;
  assign n24773 = n8418 & n22362;
  assign n24774 = n8860 & n22359;
  assign n24775 = ~n24773 & ~n24774;
  assign n24776 = ~n24772 & n24775;
  assign n24777 = ~n8421 & n24776;
  assign n24778 = n23345 & n24776;
  assign n24779 = ~n24777 & ~n24778;
  assign n24780 =  a[8]  & ~n24779;
  assign n24781 = ~ a[8]  & n24779;
  assign n24782 = ~n24780 & ~n24781;
  assign n24783 = n24771 & ~n24782;
  assign n24784 = n24359 & n24551;
  assign n24785 = ~n24552 & ~n24784;
  assign n24786 = n9331 & n22359;
  assign n24787 = n8418 & n22365;
  assign n24788 = n8860 & n22362;
  assign n24789 = ~n24787 & ~n24788;
  assign n24790 = ~n24786 & n24789;
  assign n24791 = ~n8421 & n24790;
  assign n24792 = ~n23368 & n24790;
  assign n24793 = ~n24791 & ~n24792;
  assign n24794 =  a[8]  & ~n24793;
  assign n24795 = ~ a[8]  & n24793;
  assign n24796 = ~n24794 & ~n24795;
  assign n24797 = n24785 & ~n24796;
  assign n24798 = n24377 & n24549;
  assign n24799 = ~n24550 & ~n24798;
  assign n24800 = n9331 & n22362;
  assign n24801 = n8418 & n22368;
  assign n24802 = n8860 & n22365;
  assign n24803 = ~n24801 & ~n24802;
  assign n24804 = ~n24800 & n24803;
  assign n24805 = ~n8421 & n24804;
  assign n24806 = n23320 & n24804;
  assign n24807 = ~n24805 & ~n24806;
  assign n24808 =  a[8]  & ~n24807;
  assign n24809 = ~ a[8]  & n24807;
  assign n24810 = ~n24808 & ~n24809;
  assign n24811 = n24799 & ~n24810;
  assign n24812 = n9331 & n22365;
  assign n24813 = n8418 & n22371;
  assign n24814 = n8860 & n22368;
  assign n24815 = ~n24813 & ~n24814;
  assign n24816 = ~n24812 & n24815;
  assign n24817 = n8421 & ~n22993;
  assign n24818 = n24816 & ~n24817;
  assign n24819 =  a[8]  & ~n24818;
  assign n24820 = ~n24818 & ~n24819;
  assign n24821 =  a[8]  & ~n24819;
  assign n24822 = ~n24820 & ~n24821;
  assign n24823 = n24545 & ~n24547;
  assign n24824 = ~n24548 & ~n24823;
  assign n24825 = ~n24822 & n24824;
  assign n24826 = ~n24822 & ~n24825;
  assign n24827 = n24824 & ~n24825;
  assign n24828 = ~n24826 & ~n24827;
  assign n24829 = n9331 & n22368;
  assign n24830 = n8418 & n22374;
  assign n24831 = n8860 & n22371;
  assign n24832 = ~n24830 & ~n24831;
  assign n24833 = ~n24829 & n24832;
  assign n24834 = n8421 & n23006;
  assign n24835 = n24833 & ~n24834;
  assign n24836 =  a[8]  & ~n24835;
  assign n24837 = ~n24835 & ~n24836;
  assign n24838 =  a[8]  & ~n24836;
  assign n24839 = ~n24837 & ~n24838;
  assign n24840 = ~n24540 & ~n24544;
  assign n24841 = ~n24543 & ~n24544;
  assign n24842 = ~n24840 & ~n24841;
  assign n24843 = ~n24839 & ~n24842;
  assign n24844 = ~n24839 & ~n24843;
  assign n24845 = ~n24842 & ~n24843;
  assign n24846 = ~n24844 & ~n24845;
  assign n24847 = n9331 & n22371;
  assign n24848 = n8418 & n22377;
  assign n24849 = n8860 & n22374;
  assign n24850 = ~n24848 & ~n24849;
  assign n24851 = ~n24847 & n24850;
  assign n24852 = n8421 & n23025;
  assign n24853 = n24851 & ~n24852;
  assign n24854 =  a[8]  & ~n24853;
  assign n24855 = ~n24853 & ~n24854;
  assign n24856 =  a[8]  & ~n24854;
  assign n24857 = ~n24855 & ~n24856;
  assign n24858 = ~n24535 & ~n24539;
  assign n24859 = ~n24538 & ~n24539;
  assign n24860 = ~n24858 & ~n24859;
  assign n24861 = ~n24857 & ~n24860;
  assign n24862 = ~n24857 & ~n24861;
  assign n24863 = ~n24860 & ~n24861;
  assign n24864 = ~n24862 & ~n24863;
  assign n24865 = n24436 & n24533;
  assign n24866 = ~n24534 & ~n24865;
  assign n24867 = n9331 & n22374;
  assign n24868 = n8418 & n22380;
  assign n24869 = n8860 & n22377;
  assign n24870 = ~n24868 & ~n24869;
  assign n24871 = ~n24867 & n24870;
  assign n24872 = ~n8421 & n24871;
  assign n24873 = ~n22569 & n24871;
  assign n24874 = ~n24872 & ~n24873;
  assign n24875 =  a[8]  & ~n24874;
  assign n24876 = ~ a[8]  & n24874;
  assign n24877 = ~n24875 & ~n24876;
  assign n24878 = n24866 & ~n24877;
  assign n24879 = n24529 & ~n24531;
  assign n24880 = ~n24532 & ~n24879;
  assign n24881 = n9331 & n22377;
  assign n24882 = n8418 & n22384;
  assign n24883 = n8860 & n22380;
  assign n24884 = ~n24882 & ~n24883;
  assign n24885 = ~n24881 & n24884;
  assign n24886 = ~n8421 & n24885;
  assign n24887 = n22834 & n24885;
  assign n24888 = ~n24886 & ~n24887;
  assign n24889 =  a[8]  & ~n24888;
  assign n24890 = ~ a[8]  & n24888;
  assign n24891 = ~n24889 & ~n24890;
  assign n24892 = n24880 & ~n24891;
  assign n24893 = n24468 & n24527;
  assign n24894 = ~n24528 & ~n24893;
  assign n24895 = n9331 & n22380;
  assign n24896 = n8418 & n22387;
  assign n24897 = n8860 & n22384;
  assign n24898 = ~n24896 & ~n24897;
  assign n24899 = ~n24895 & n24898;
  assign n24900 = ~n8421 & n24899;
  assign n24901 = ~n22850 & n24899;
  assign n24902 = ~n24900 & ~n24901;
  assign n24903 =  a[8]  & ~n24902;
  assign n24904 = ~ a[8]  & n24902;
  assign n24905 = ~n24903 & ~n24904;
  assign n24906 = n24894 & ~n24905;
  assign n24907 = n9331 & n22384;
  assign n24908 = n8418 & n22390;
  assign n24909 = n8860 & n22387;
  assign n24910 = ~n24908 & ~n24909;
  assign n24911 = ~n24907 & n24910;
  assign n24912 = n8421 & n22806;
  assign n24913 = n24911 & ~n24912;
  assign n24914 =  a[8]  & ~n24913;
  assign n24915 = ~n24913 & ~n24914;
  assign n24916 =  a[8]  & ~n24914;
  assign n24917 = ~n24915 & ~n24916;
  assign n24918 = n24523 & ~n24525;
  assign n24919 = ~n24526 & ~n24918;
  assign n24920 = ~n24917 & n24919;
  assign n24921 = ~n24917 & ~n24920;
  assign n24922 = n24919 & ~n24920;
  assign n24923 = ~n24921 & ~n24922;
  assign n24924 = ~n24510 & ~n24522;
  assign n24925 = ~n24521 & ~n24522;
  assign n24926 = ~n24924 & ~n24925;
  assign n24927 = n9331 & n22387;
  assign n24928 = n8418 & n22393;
  assign n24929 = n8860 & n22390;
  assign n24930 = ~n24928 & ~n24929;
  assign n24931 = ~n24927 & n24930;
  assign n24932 = ~n8421 & n24931;
  assign n24933 = ~n22582 & n24931;
  assign n24934 = ~n24932 & ~n24933;
  assign n24935 =  a[8]  & ~n24934;
  assign n24936 = ~ a[8]  & n24934;
  assign n24937 = ~n24935 & ~n24936;
  assign n24938 = ~n24926 & ~n24937;
  assign n24939 = n9331 & n22390;
  assign n24940 = n8418 & n22396;
  assign n24941 = n8860 & n22393;
  assign n24942 = ~n24940 & ~n24941;
  assign n24943 = ~n24939 & n24942;
  assign n24944 = n8421 & n22649;
  assign n24945 = n24943 & ~n24944;
  assign n24946 =  a[8]  & ~n24945;
  assign n24947 = ~n24945 & ~n24946;
  assign n24948 =  a[8]  & ~n24946;
  assign n24949 = ~n24947 & ~n24948;
  assign n24950 = ~n24494 & n24505;
  assign n24951 = ~n24506 & ~n24950;
  assign n24952 = ~n24949 & n24951;
  assign n24953 = ~n24949 & ~n24952;
  assign n24954 = n24951 & ~n24952;
  assign n24955 = ~n24953 & ~n24954;
  assign n24956 = n24491 & ~n24493;
  assign n24957 = ~n24494 & ~n24956;
  assign n24958 = n9331 & n22393;
  assign n24959 = n8418 & n22399;
  assign n24960 = n8860 & n22396;
  assign n24961 = ~n24959 & ~n24960;
  assign n24962 = ~n24958 & n24961;
  assign n24963 = ~n8421 & n24962;
  assign n24964 = ~n22671 & n24962;
  assign n24965 = ~n24963 & ~n24964;
  assign n24966 =  a[8]  & ~n24965;
  assign n24967 = ~ a[8]  & n24965;
  assign n24968 = ~n24966 & ~n24967;
  assign n24969 = n24957 & ~n24968;
  assign n24970 = n8860 & ~n22406;
  assign n24971 = n9331 & n22402;
  assign n24972 = ~n24970 & ~n24971;
  assign n24973 = n8421 & ~n22609;
  assign n24974 = n24972 & ~n24973;
  assign n24975 =  a[8]  & ~n24974;
  assign n24976 =  a[8]  & ~n24975;
  assign n24977 = ~n24974 & ~n24975;
  assign n24978 = ~n24976 & ~n24977;
  assign n24979 = ~n8416 & ~n22406;
  assign n24980 =  a[8]  & ~n24979;
  assign n24981 = ~n24978 & n24980;
  assign n24982 = n9331 & n22399;
  assign n24983 = n8418 & ~n22406;
  assign n24984 = n8860 & n22402;
  assign n24985 = ~n24983 & ~n24984;
  assign n24986 = ~n24982 & n24985;
  assign n24987 = ~n8421 & n24986;
  assign n24988 = n22625 & n24986;
  assign n24989 = ~n24987 & ~n24988;
  assign n24990 =  a[8]  & ~n24989;
  assign n24991 = ~ a[8]  & n24989;
  assign n24992 = ~n24990 & ~n24991;
  assign n24993 = n24981 & ~n24992;
  assign n24994 = n24492 & n24993;
  assign n24995 = n24993 & ~n24994;
  assign n24996 = n24492 & ~n24994;
  assign n24997 = ~n24995 & ~n24996;
  assign n24998 = n9331 & n22396;
  assign n24999 = n8418 & n22402;
  assign n25000 = n8860 & n22399;
  assign n25001 = ~n24999 & ~n25000;
  assign n25002 = ~n24998 & n25001;
  assign n25003 = n8421 & n22595;
  assign n25004 = n25002 & ~n25003;
  assign n25005 =  a[8]  & ~n25004;
  assign n25006 =  a[8]  & ~n25005;
  assign n25007 = ~n25004 & ~n25005;
  assign n25008 = ~n25006 & ~n25007;
  assign n25009 = ~n24997 & ~n25008;
  assign n25010 = ~n24994 & ~n25009;
  assign n25011 = ~n24957 & n24968;
  assign n25012 = ~n24969 & ~n25011;
  assign n25013 = ~n25010 & n25012;
  assign n25014 = ~n24969 & ~n25013;
  assign n25015 = ~n24955 & ~n25014;
  assign n25016 = ~n24952 & ~n25015;
  assign n25017 = n24926 & n24937;
  assign n25018 = ~n24938 & ~n25017;
  assign n25019 = ~n25016 & n25018;
  assign n25020 = ~n24938 & ~n25019;
  assign n25021 = ~n24923 & ~n25020;
  assign n25022 = ~n24920 & ~n25021;
  assign n25023 = n24894 & ~n24906;
  assign n25024 = ~n24905 & ~n24906;
  assign n25025 = ~n25023 & ~n25024;
  assign n25026 = ~n25022 & ~n25025;
  assign n25027 = ~n24906 & ~n25026;
  assign n25028 = n24880 & ~n24892;
  assign n25029 = ~n24891 & ~n24892;
  assign n25030 = ~n25028 & ~n25029;
  assign n25031 = ~n25027 & ~n25030;
  assign n25032 = ~n24892 & ~n25031;
  assign n25033 = ~n24866 & n24877;
  assign n25034 = ~n24878 & ~n25033;
  assign n25035 = ~n25032 & n25034;
  assign n25036 = ~n24878 & ~n25035;
  assign n25037 = ~n24864 & ~n25036;
  assign n25038 = ~n24861 & ~n25037;
  assign n25039 = ~n24846 & ~n25038;
  assign n25040 = ~n24843 & ~n25039;
  assign n25041 = ~n24828 & ~n25040;
  assign n25042 = ~n24825 & ~n25041;
  assign n25043 = n24799 & ~n24811;
  assign n25044 = ~n24810 & ~n24811;
  assign n25045 = ~n25043 & ~n25044;
  assign n25046 = ~n25042 & ~n25045;
  assign n25047 = ~n24811 & ~n25046;
  assign n25048 = n24785 & ~n24797;
  assign n25049 = ~n24796 & ~n24797;
  assign n25050 = ~n25048 & ~n25049;
  assign n25051 = ~n25047 & ~n25050;
  assign n25052 = ~n24797 & ~n25051;
  assign n25053 = ~n24771 & n24782;
  assign n25054 = ~n24783 & ~n25053;
  assign n25055 = ~n25052 & n25054;
  assign n25056 = ~n24783 & ~n25055;
  assign n25057 = ~n24769 & ~n25056;
  assign n25058 = ~n24766 & ~n25057;
  assign n25059 = ~n24751 & ~n25058;
  assign n25060 = ~n24748 & ~n25059;
  assign n25061 = ~n24733 & ~n25060;
  assign n25062 = ~n24730 & ~n25061;
  assign n25063 = n24704 & ~n24716;
  assign n25064 = ~n24715 & ~n24716;
  assign n25065 = ~n25063 & ~n25064;
  assign n25066 = ~n25062 & ~n25065;
  assign n25067 = ~n24716 & ~n25066;
  assign n25068 = n24690 & ~n24702;
  assign n25069 = ~n24701 & ~n24702;
  assign n25070 = ~n25068 & ~n25069;
  assign n25071 = ~n25067 & ~n25070;
  assign n25072 = ~n24702 & ~n25071;
  assign n25073 = ~n24676 & n24687;
  assign n25074 = ~n24688 & ~n25073;
  assign n25075 = ~n25072 & n25074;
  assign n25076 = ~n24688 & ~n25075;
  assign n25077 = ~n24674 & ~n25076;
  assign n25078 = ~n24671 & ~n25077;
  assign n25079 = ~n24656 & ~n25078;
  assign n25080 = ~n24653 & ~n25079;
  assign n25081 = n24624 & ~n24639;
  assign n25082 = ~n24638 & ~n24639;
  assign n25083 = ~n25081 & ~n25082;
  assign n25084 = ~n25080 & ~n25083;
  assign n25085 = ~n24639 & ~n25084;
  assign n25086 = n24607 & ~n24622;
  assign n25087 = ~n24621 & ~n24622;
  assign n25088 = ~n25086 & ~n25087;
  assign n25089 = ~n25085 & ~n25088;
  assign n25090 = ~n24622 & ~n25089;
  assign n25091 = n24591 & ~n24605;
  assign n25092 = ~n24604 & ~n24605;
  assign n25093 = ~n25091 & ~n25092;
  assign n25094 = ~n25090 & ~n25093;
  assign n25095 = ~n24605 & ~n25094;
  assign n25096 = n7983 & n22329;
  assign n25097 = n7291 & n22335;
  assign n25098 = n7632 & n22332;
  assign n25099 = ~n25097 & ~n25098;
  assign n25100 = ~n25096 & n25099;
  assign n25101 = n7294 & ~n24633;
  assign n25102 = n25100 & ~n25101;
  assign n25103 =  a[11]  & ~n25102;
  assign n25104 = ~n25102 & ~n25103;
  assign n25105 =  a[11]  & ~n25103;
  assign n25106 = ~n25104 & ~n25105;
  assign n25107 = ~n24148 & ~n24152;
  assign n25108 = n6233 & n22347;
  assign n25109 = n5663 & n22353;
  assign n25110 = n5939 & n22350;
  assign n25111 = ~n25109 & ~n25110;
  assign n25112 = ~n25108 & n25111;
  assign n25113 = n5666 & ~n23659;
  assign n25114 = n25112 & ~n25113;
  assign n25115 =  a[17]  & ~n25114;
  assign n25116 = ~n25114 & ~n25115;
  assign n25117 =  a[17]  & ~n25115;
  assign n25118 = ~n25116 & ~n25117;
  assign n25119 = ~n24119 & ~n24123;
  assign n25120 = n4694 & n22365;
  assign n25121 = n4533 & n22371;
  assign n25122 = n4604 & n22368;
  assign n25123 = ~n25121 & ~n25122;
  assign n25124 = ~n25120 & n25123;
  assign n25125 = n4536 & ~n22993;
  assign n25126 = n25124 & ~n25125;
  assign n25127 =  a[23]  & ~n25126;
  assign n25128 = ~n25126 & ~n25127;
  assign n25129 =  a[23]  & ~n25127;
  assign n25130 = ~n25128 & ~n25129;
  assign n25131 = ~n24092 & ~n24096;
  assign n25132 = n3457 & n22384;
  assign n25133 = n3542 & n22390;
  assign n25134 = n3606 & n22387;
  assign n25135 = ~n25133 & ~n25134;
  assign n25136 = ~n25132 & n25135;
  assign n25137 = n3368 & n22806;
  assign n25138 = n25136 & ~n25137;
  assign n25139 =  a[29]  & ~n25138;
  assign n25140 = ~n25138 & ~n25139;
  assign n25141 =  a[29]  & ~n25139;
  assign n25142 = ~n25140 & ~n25141;
  assign n25143 = ~n24065 & ~n24069;
  assign n25144 = n1611 & n5748;
  assign n25145 = n4269 & n25144;
  assign n25146 = n691 & n25145;
  assign n25147 = n204 & n25146;
  assign n25148 = n13560 & n25147;
  assign n25149 = n12932 & n25148;
  assign n25150 = n12909 & n25149;
  assign n25151 = n15924 & n25150;
  assign n25152 = n515 & n25151;
  assign n25153 = ~n278 & n25152;
  assign n25154 = ~n135 & n25153;
  assign n25155 = ~n568 & n25154;
  assign n25156 = ~n331 & n25155;
  assign n25157 = ~n225 & n25156;
  assign n25158 = n3020 & n22393;
  assign n25159 = n3028 & n22396;
  assign n25160 = n3023 & n22399;
  assign n25161 = n75 & n22671;
  assign n25162 = ~n25160 & ~n25161;
  assign n25163 = ~n25159 & n25162;
  assign n25164 = ~n25158 & n25163;
  assign n25165 = ~n25157 & ~n25164;
  assign n25166 = ~n25157 & ~n25165;
  assign n25167 = ~n25164 & ~n25165;
  assign n25168 = ~n25166 & ~n25167;
  assign n25169 = ~n25143 & ~n25168;
  assign n25170 = ~n25143 & ~n25169;
  assign n25171 = ~n25168 & ~n25169;
  assign n25172 = ~n25170 & ~n25171;
  assign n25173 = ~n25142 & ~n25172;
  assign n25174 = ~n25142 & ~n25173;
  assign n25175 = ~n25172 & ~n25173;
  assign n25176 = ~n25174 & ~n25175;
  assign n25177 = ~n24073 & ~n24079;
  assign n25178 = n25176 & n25177;
  assign n25179 = ~n25176 & ~n25177;
  assign n25180 = ~n25178 & ~n25179;
  assign n25181 = n3884 & n22374;
  assign n25182 = n3967 & n22380;
  assign n25183 = n4046 & n22377;
  assign n25184 = ~n25182 & ~n25183;
  assign n25185 = ~n25181 & n25184;
  assign n25186 = ~n4050 & n25185;
  assign n25187 = ~n22569 & n25185;
  assign n25188 = ~n25186 & ~n25187;
  assign n25189 =  a[26]  & ~n25188;
  assign n25190 = ~ a[26]  & n25188;
  assign n25191 = ~n25189 & ~n25190;
  assign n25192 = n25180 & ~n25191;
  assign n25193 = n25180 & ~n25192;
  assign n25194 = ~n25191 & ~n25192;
  assign n25195 = ~n25193 & ~n25194;
  assign n25196 = ~n25131 & ~n25195;
  assign n25197 = ~n25131 & ~n25196;
  assign n25198 = ~n25195 & ~n25196;
  assign n25199 = ~n25197 & ~n25198;
  assign n25200 = ~n25130 & ~n25199;
  assign n25201 = ~n25130 & ~n25200;
  assign n25202 = ~n25199 & ~n25200;
  assign n25203 = ~n25201 & ~n25202;
  assign n25204 = ~n24100 & ~n24106;
  assign n25205 = n25203 & n25204;
  assign n25206 = ~n25203 & ~n25204;
  assign n25207 = ~n25205 & ~n25206;
  assign n25208 = n5496 & n22356;
  assign n25209 = n4935 & n22362;
  assign n25210 = n5407 & n22359;
  assign n25211 = ~n25209 & ~n25210;
  assign n25212 = ~n25208 & n25211;
  assign n25213 = ~n4938 & n25212;
  assign n25214 = n23345 & n25212;
  assign n25215 = ~n25213 & ~n25214;
  assign n25216 =  a[20]  & ~n25215;
  assign n25217 = ~ a[20]  & n25215;
  assign n25218 = ~n25216 & ~n25217;
  assign n25219 = n25207 & ~n25218;
  assign n25220 = n25207 & ~n25219;
  assign n25221 = ~n25218 & ~n25219;
  assign n25222 = ~n25220 & ~n25221;
  assign n25223 = ~n25119 & ~n25222;
  assign n25224 = ~n25119 & ~n25223;
  assign n25225 = ~n25222 & ~n25223;
  assign n25226 = ~n25224 & ~n25225;
  assign n25227 = ~n25118 & ~n25226;
  assign n25228 = ~n25118 & ~n25227;
  assign n25229 = ~n25226 & ~n25227;
  assign n25230 = ~n25228 & ~n25229;
  assign n25231 = ~n24127 & ~n24133;
  assign n25232 = n25230 & n25231;
  assign n25233 = ~n25230 & ~n25231;
  assign n25234 = ~n25232 & ~n25233;
  assign n25235 = n7101 & n22338;
  assign n25236 = n6402 & n22344;
  assign n25237 = n6951 & n22341;
  assign n25238 = ~n25236 & ~n25237;
  assign n25239 = ~n25235 & n25238;
  assign n25240 = ~n6397 & n25239;
  assign n25241 = n24188 & n25239;
  assign n25242 = ~n25240 & ~n25241;
  assign n25243 =  a[14]  & ~n25242;
  assign n25244 = ~ a[14]  & n25242;
  assign n25245 = ~n25243 & ~n25244;
  assign n25246 = n25234 & ~n25245;
  assign n25247 = n25234 & ~n25246;
  assign n25248 = ~n25245 & ~n25246;
  assign n25249 = ~n25247 & ~n25248;
  assign n25250 = ~n25107 & ~n25249;
  assign n25251 = ~n25107 & ~n25250;
  assign n25252 = ~n25249 & ~n25250;
  assign n25253 = ~n25251 & ~n25252;
  assign n25254 = ~n25106 & ~n25253;
  assign n25255 = ~n25106 & ~n25254;
  assign n25256 = ~n25253 & ~n25254;
  assign n25257 = ~n25255 & ~n25256;
  assign n25258 = ~n24156 & ~n24590;
  assign n25259 = n25257 & n25258;
  assign n25260 = ~n25257 & ~n25258;
  assign n25261 = ~n25259 & ~n25260;
  assign n25262 = n9331 & n22320;
  assign n25263 = n8418 & n22326;
  assign n25264 = n8860 & n22323;
  assign n25265 = ~n25263 & ~n25264;
  assign n25266 = ~n25262 & n25265;
  assign n25267 = ~n8421 & n25266;
  assign n25268 = ~n22508 & ~n22511;
  assign n25269 = ~n22509 & n22512;
  assign n25270 = ~n25268 & ~n25269;
  assign n25271 = n25266 & n25270;
  assign n25272 = ~n25267 & ~n25271;
  assign n25273 =  a[8]  & ~n25272;
  assign n25274 = ~ a[8]  & n25272;
  assign n25275 = ~n25273 & ~n25274;
  assign n25276 = n25261 & ~n25275;
  assign n25277 = n25261 & ~n25276;
  assign n25278 = ~n25275 & ~n25276;
  assign n25279 = ~n25277 & ~n25278;
  assign n25280 = ~n25095 & ~n25279;
  assign n25281 = ~n25095 & ~n25280;
  assign n25282 = ~n25279 & ~n25280;
  assign n25283 = ~n25281 & ~n25282;
  assign n25284 = ~n22535 & ~n25283;
  assign n25285 = ~n22535 & ~n25284;
  assign n25286 = ~n25283 & ~n25284;
  assign n25287 = ~n25285 & ~n25286;
  assign n25288 = n71 & n22315;
  assign n25289 = n9867 & n22320;
  assign n25290 = n10434 & n22312;
  assign n25291 = ~n25289 & ~n25290;
  assign n25292 = ~n25288 & n25291;
  assign n25293 = n22516 & ~n22519;
  assign n25294 = ~n22520 & ~n25293;
  assign n25295 = n9870 & n25294;
  assign n25296 = n25292 & ~n25295;
  assign n25297 =  a[5]  & ~n25296;
  assign n25298 = ~n25296 & ~n25297;
  assign n25299 =  a[5]  & ~n25297;
  assign n25300 = ~n25298 & ~n25299;
  assign n25301 = ~n25090 & ~n25094;
  assign n25302 = ~n25093 & ~n25094;
  assign n25303 = ~n25301 & ~n25302;
  assign n25304 = ~n25300 & ~n25303;
  assign n25305 = ~n25300 & ~n25304;
  assign n25306 = ~n25303 & ~n25304;
  assign n25307 = ~n25305 & ~n25306;
  assign n25308 = n71 & n22312;
  assign n25309 = n9867 & n22323;
  assign n25310 = n10434 & n22320;
  assign n25311 = ~n25309 & ~n25310;
  assign n25312 = ~n25308 & n25311;
  assign n25313 = ~n22512 & ~n22515;
  assign n25314 = ~n22513 & n22516;
  assign n25315 = ~n25313 & ~n25314;
  assign n25316 = n9870 & ~n25315;
  assign n25317 = n25312 & ~n25316;
  assign n25318 =  a[5]  & ~n25317;
  assign n25319 = ~n25317 & ~n25318;
  assign n25320 =  a[5]  & ~n25318;
  assign n25321 = ~n25319 & ~n25320;
  assign n25322 = ~n25085 & ~n25089;
  assign n25323 = ~n25088 & ~n25089;
  assign n25324 = ~n25322 & ~n25323;
  assign n25325 = ~n25321 & ~n25324;
  assign n25326 = ~n25321 & ~n25325;
  assign n25327 = ~n25324 & ~n25325;
  assign n25328 = ~n25326 & ~n25327;
  assign n25329 = n71 & n22320;
  assign n25330 = n9867 & n22326;
  assign n25331 = n10434 & n22323;
  assign n25332 = ~n25330 & ~n25331;
  assign n25333 = ~n25329 & n25332;
  assign n25334 = n9870 & ~n25270;
  assign n25335 = n25333 & ~n25334;
  assign n25336 =  a[5]  & ~n25335;
  assign n25337 = ~n25335 & ~n25336;
  assign n25338 =  a[5]  & ~n25336;
  assign n25339 = ~n25337 & ~n25338;
  assign n25340 = ~n25080 & ~n25084;
  assign n25341 = ~n25083 & ~n25084;
  assign n25342 = ~n25340 & ~n25341;
  assign n25343 = ~n25339 & ~n25342;
  assign n25344 = ~n25339 & ~n25343;
  assign n25345 = ~n25342 & ~n25343;
  assign n25346 = ~n25344 & ~n25345;
  assign n25347 = n24656 & n25078;
  assign n25348 = ~n25079 & ~n25347;
  assign n25349 = n71 & n22323;
  assign n25350 = n9867 & n22329;
  assign n25351 = n10434 & n22326;
  assign n25352 = ~n25350 & ~n25351;
  assign n25353 = ~n25349 & n25352;
  assign n25354 = ~n9870 & n25353;
  assign n25355 = ~n24599 & n25353;
  assign n25356 = ~n25354 & ~n25355;
  assign n25357 =  a[5]  & ~n25356;
  assign n25358 = ~ a[5]  & n25356;
  assign n25359 = ~n25357 & ~n25358;
  assign n25360 = n25348 & ~n25359;
  assign n25361 = n24674 & n25076;
  assign n25362 = ~n25077 & ~n25361;
  assign n25363 = n71 & n22326;
  assign n25364 = n9867 & n22332;
  assign n25365 = n10434 & n22329;
  assign n25366 = ~n25364 & ~n25365;
  assign n25367 = ~n25363 & n25366;
  assign n25368 = ~n9870 & n25367;
  assign n25369 = n24616 & n25367;
  assign n25370 = ~n25368 & ~n25369;
  assign n25371 =  a[5]  & ~n25370;
  assign n25372 = ~ a[5]  & n25370;
  assign n25373 = ~n25371 & ~n25372;
  assign n25374 = n25362 & ~n25373;
  assign n25375 = n71 & n22329;
  assign n25376 = n9867 & n22335;
  assign n25377 = n10434 & n22332;
  assign n25378 = ~n25376 & ~n25377;
  assign n25379 = ~n25375 & n25378;
  assign n25380 = n9870 & ~n24633;
  assign n25381 = n25379 & ~n25380;
  assign n25382 =  a[5]  & ~n25381;
  assign n25383 = ~n25381 & ~n25382;
  assign n25384 =  a[5]  & ~n25382;
  assign n25385 = ~n25383 & ~n25384;
  assign n25386 = n25072 & ~n25074;
  assign n25387 = ~n25075 & ~n25386;
  assign n25388 = ~n25385 & n25387;
  assign n25389 = ~n25385 & ~n25388;
  assign n25390 = n25387 & ~n25388;
  assign n25391 = ~n25389 & ~n25390;
  assign n25392 = n71 & n22332;
  assign n25393 = n9867 & n22338;
  assign n25394 = n10434 & n22335;
  assign n25395 = ~n25393 & ~n25394;
  assign n25396 = ~n25392 & n25395;
  assign n25397 = n9870 & n22542;
  assign n25398 = n25396 & ~n25397;
  assign n25399 =  a[5]  & ~n25398;
  assign n25400 = ~n25398 & ~n25399;
  assign n25401 =  a[5]  & ~n25399;
  assign n25402 = ~n25400 & ~n25401;
  assign n25403 = ~n25067 & ~n25071;
  assign n25404 = ~n25070 & ~n25071;
  assign n25405 = ~n25403 & ~n25404;
  assign n25406 = ~n25402 & ~n25405;
  assign n25407 = ~n25402 & ~n25406;
  assign n25408 = ~n25405 & ~n25406;
  assign n25409 = ~n25407 & ~n25408;
  assign n25410 = n71 & n22335;
  assign n25411 = n9867 & n22341;
  assign n25412 = n10434 & n22338;
  assign n25413 = ~n25411 & ~n25412;
  assign n25414 = ~n25410 & n25413;
  assign n25415 = n9870 & ~n24167;
  assign n25416 = n25414 & ~n25415;
  assign n25417 =  a[5]  & ~n25416;
  assign n25418 = ~n25416 & ~n25417;
  assign n25419 =  a[5]  & ~n25417;
  assign n25420 = ~n25418 & ~n25419;
  assign n25421 = ~n25062 & ~n25066;
  assign n25422 = ~n25065 & ~n25066;
  assign n25423 = ~n25421 & ~n25422;
  assign n25424 = ~n25420 & ~n25423;
  assign n25425 = ~n25420 & ~n25424;
  assign n25426 = ~n25423 & ~n25424;
  assign n25427 = ~n25425 & ~n25426;
  assign n25428 = n24733 & n25060;
  assign n25429 = ~n25061 & ~n25428;
  assign n25430 = n71 & n22338;
  assign n25431 = n9867 & n22344;
  assign n25432 = n10434 & n22341;
  assign n25433 = ~n25431 & ~n25432;
  assign n25434 = ~n25430 & n25433;
  assign n25435 = ~n9870 & n25434;
  assign n25436 = n24188 & n25434;
  assign n25437 = ~n25435 & ~n25436;
  assign n25438 =  a[5]  & ~n25437;
  assign n25439 = ~ a[5]  & n25437;
  assign n25440 = ~n25438 & ~n25439;
  assign n25441 = n25429 & ~n25440;
  assign n25442 = n24751 & n25058;
  assign n25443 = ~n25059 & ~n25442;
  assign n25444 = n71 & n22341;
  assign n25445 = n9867 & n22347;
  assign n25446 = n10434 & n22344;
  assign n25447 = ~n25445 & ~n25446;
  assign n25448 = ~n25444 & n25447;
  assign n25449 = ~n9870 & n25448;
  assign n25450 = ~n24142 & n25448;
  assign n25451 = ~n25449 & ~n25450;
  assign n25452 =  a[5]  & ~n25451;
  assign n25453 = ~ a[5]  & n25451;
  assign n25454 = ~n25452 & ~n25453;
  assign n25455 = n25443 & ~n25454;
  assign n25456 = n24769 & n25056;
  assign n25457 = ~n25057 & ~n25456;
  assign n25458 = n71 & n22344;
  assign n25459 = n9867 & n22350;
  assign n25460 = n10434 & n22347;
  assign n25461 = ~n25459 & ~n25460;
  assign n25462 = ~n25458 & n25461;
  assign n25463 = ~n9870 & n25462;
  assign n25464 = n23642 & n25462;
  assign n25465 = ~n25463 & ~n25464;
  assign n25466 =  a[5]  & ~n25465;
  assign n25467 = ~ a[5]  & n25465;
  assign n25468 = ~n25466 & ~n25467;
  assign n25469 = n25457 & ~n25468;
  assign n25470 = n71 & n22347;
  assign n25471 = n9867 & n22353;
  assign n25472 = n10434 & n22350;
  assign n25473 = ~n25471 & ~n25472;
  assign n25474 = ~n25470 & n25473;
  assign n25475 = n9870 & ~n23659;
  assign n25476 = n25474 & ~n25475;
  assign n25477 =  a[5]  & ~n25476;
  assign n25478 = ~n25476 & ~n25477;
  assign n25479 =  a[5]  & ~n25477;
  assign n25480 = ~n25478 & ~n25479;
  assign n25481 = n25052 & ~n25054;
  assign n25482 = ~n25055 & ~n25481;
  assign n25483 = ~n25480 & n25482;
  assign n25484 = ~n25480 & ~n25483;
  assign n25485 = n25482 & ~n25483;
  assign n25486 = ~n25484 & ~n25485;
  assign n25487 = n71 & n22350;
  assign n25488 = n9867 & n22356;
  assign n25489 = n10434 & n22353;
  assign n25490 = ~n25488 & ~n25489;
  assign n25491 = ~n25487 & n25490;
  assign n25492 = n9870 & n23672;
  assign n25493 = n25491 & ~n25492;
  assign n25494 =  a[5]  & ~n25493;
  assign n25495 = ~n25493 & ~n25494;
  assign n25496 =  a[5]  & ~n25494;
  assign n25497 = ~n25495 & ~n25496;
  assign n25498 = ~n25047 & ~n25051;
  assign n25499 = ~n25050 & ~n25051;
  assign n25500 = ~n25498 & ~n25499;
  assign n25501 = ~n25497 & ~n25500;
  assign n25502 = ~n25497 & ~n25501;
  assign n25503 = ~n25500 & ~n25501;
  assign n25504 = ~n25502 & ~n25503;
  assign n25505 = n71 & n22353;
  assign n25506 = n9867 & n22359;
  assign n25507 = n10434 & n22356;
  assign n25508 = ~n25506 & ~n25507;
  assign n25509 = ~n25505 & n25508;
  assign n25510 = n9870 & ~n22556;
  assign n25511 = n25509 & ~n25510;
  assign n25512 =  a[5]  & ~n25511;
  assign n25513 = ~n25511 & ~n25512;
  assign n25514 =  a[5]  & ~n25512;
  assign n25515 = ~n25513 & ~n25514;
  assign n25516 = ~n25042 & ~n25046;
  assign n25517 = ~n25045 & ~n25046;
  assign n25518 = ~n25516 & ~n25517;
  assign n25519 = ~n25515 & ~n25518;
  assign n25520 = ~n25515 & ~n25519;
  assign n25521 = ~n25518 & ~n25519;
  assign n25522 = ~n25520 & ~n25521;
  assign n25523 = n24828 & n25040;
  assign n25524 = ~n25041 & ~n25523;
  assign n25525 = n71 & n22356;
  assign n25526 = n9867 & n22362;
  assign n25527 = n10434 & n22359;
  assign n25528 = ~n25526 & ~n25527;
  assign n25529 = ~n25525 & n25528;
  assign n25530 = ~n9870 & n25529;
  assign n25531 = n23345 & n25529;
  assign n25532 = ~n25530 & ~n25531;
  assign n25533 =  a[5]  & ~n25532;
  assign n25534 = ~ a[5]  & n25532;
  assign n25535 = ~n25533 & ~n25534;
  assign n25536 = n25524 & ~n25535;
  assign n25537 = n24846 & n25038;
  assign n25538 = ~n25039 & ~n25537;
  assign n25539 = n71 & n22359;
  assign n25540 = n9867 & n22365;
  assign n25541 = n10434 & n22362;
  assign n25542 = ~n25540 & ~n25541;
  assign n25543 = ~n25539 & n25542;
  assign n25544 = ~n9870 & n25543;
  assign n25545 = ~n23368 & n25543;
  assign n25546 = ~n25544 & ~n25545;
  assign n25547 =  a[5]  & ~n25546;
  assign n25548 = ~ a[5]  & n25546;
  assign n25549 = ~n25547 & ~n25548;
  assign n25550 = n25538 & ~n25549;
  assign n25551 = n24864 & n25036;
  assign n25552 = ~n25037 & ~n25551;
  assign n25553 = n71 & n22362;
  assign n25554 = n9867 & n22368;
  assign n25555 = n10434 & n22365;
  assign n25556 = ~n25554 & ~n25555;
  assign n25557 = ~n25553 & n25556;
  assign n25558 = ~n9870 & n25557;
  assign n25559 = n23320 & n25557;
  assign n25560 = ~n25558 & ~n25559;
  assign n25561 =  a[5]  & ~n25560;
  assign n25562 = ~ a[5]  & n25560;
  assign n25563 = ~n25561 & ~n25562;
  assign n25564 = n25552 & ~n25563;
  assign n25565 = n71 & n22365;
  assign n25566 = n9867 & n22371;
  assign n25567 = n10434 & n22368;
  assign n25568 = ~n25566 & ~n25567;
  assign n25569 = ~n25565 & n25568;
  assign n25570 = n9870 & ~n22993;
  assign n25571 = n25569 & ~n25570;
  assign n25572 =  a[5]  & ~n25571;
  assign n25573 = ~n25571 & ~n25572;
  assign n25574 =  a[5]  & ~n25572;
  assign n25575 = ~n25573 & ~n25574;
  assign n25576 = n25032 & ~n25034;
  assign n25577 = ~n25035 & ~n25576;
  assign n25578 = ~n25575 & n25577;
  assign n25579 = ~n25575 & ~n25578;
  assign n25580 = n25577 & ~n25578;
  assign n25581 = ~n25579 & ~n25580;
  assign n25582 = n71 & n22368;
  assign n25583 = n9867 & n22374;
  assign n25584 = n10434 & n22371;
  assign n25585 = ~n25583 & ~n25584;
  assign n25586 = ~n25582 & n25585;
  assign n25587 = n9870 & n23006;
  assign n25588 = n25586 & ~n25587;
  assign n25589 =  a[5]  & ~n25588;
  assign n25590 = ~n25588 & ~n25589;
  assign n25591 =  a[5]  & ~n25589;
  assign n25592 = ~n25590 & ~n25591;
  assign n25593 = ~n25027 & ~n25031;
  assign n25594 = ~n25030 & ~n25031;
  assign n25595 = ~n25593 & ~n25594;
  assign n25596 = ~n25592 & ~n25595;
  assign n25597 = ~n25592 & ~n25596;
  assign n25598 = ~n25595 & ~n25596;
  assign n25599 = ~n25597 & ~n25598;
  assign n25600 = n71 & n22371;
  assign n25601 = n9867 & n22377;
  assign n25602 = n10434 & n22374;
  assign n25603 = ~n25601 & ~n25602;
  assign n25604 = ~n25600 & n25603;
  assign n25605 = n9870 & n23025;
  assign n25606 = n25604 & ~n25605;
  assign n25607 =  a[5]  & ~n25606;
  assign n25608 = ~n25606 & ~n25607;
  assign n25609 =  a[5]  & ~n25607;
  assign n25610 = ~n25608 & ~n25609;
  assign n25611 = ~n25022 & ~n25026;
  assign n25612 = ~n25025 & ~n25026;
  assign n25613 = ~n25611 & ~n25612;
  assign n25614 = ~n25610 & ~n25613;
  assign n25615 = ~n25610 & ~n25614;
  assign n25616 = ~n25613 & ~n25614;
  assign n25617 = ~n25615 & ~n25616;
  assign n25618 = n24923 & n25020;
  assign n25619 = ~n25021 & ~n25618;
  assign n25620 = n71 & n22374;
  assign n25621 = n9867 & n22380;
  assign n25622 = n10434 & n22377;
  assign n25623 = ~n25621 & ~n25622;
  assign n25624 = ~n25620 & n25623;
  assign n25625 = ~n9870 & n25624;
  assign n25626 = ~n22569 & n25624;
  assign n25627 = ~n25625 & ~n25626;
  assign n25628 =  a[5]  & ~n25627;
  assign n25629 = ~ a[5]  & n25627;
  assign n25630 = ~n25628 & ~n25629;
  assign n25631 = n25619 & ~n25630;
  assign n25632 = n25016 & ~n25018;
  assign n25633 = ~n25019 & ~n25632;
  assign n25634 = n71 & n22377;
  assign n25635 = n9867 & n22384;
  assign n25636 = n10434 & n22380;
  assign n25637 = ~n25635 & ~n25636;
  assign n25638 = ~n25634 & n25637;
  assign n25639 = ~n9870 & n25638;
  assign n25640 = n22834 & n25638;
  assign n25641 = ~n25639 & ~n25640;
  assign n25642 =  a[5]  & ~n25641;
  assign n25643 = ~ a[5]  & n25641;
  assign n25644 = ~n25642 & ~n25643;
  assign n25645 = n25633 & ~n25644;
  assign n25646 = n24955 & n25014;
  assign n25647 = ~n25015 & ~n25646;
  assign n25648 = n71 & n22380;
  assign n25649 = n9867 & n22387;
  assign n25650 = n10434 & n22384;
  assign n25651 = ~n25649 & ~n25650;
  assign n25652 = ~n25648 & n25651;
  assign n25653 = ~n9870 & n25652;
  assign n25654 = ~n22850 & n25652;
  assign n25655 = ~n25653 & ~n25654;
  assign n25656 =  a[5]  & ~n25655;
  assign n25657 = ~ a[5]  & n25655;
  assign n25658 = ~n25656 & ~n25657;
  assign n25659 = n25647 & ~n25658;
  assign n25660 = n71 & n22384;
  assign n25661 = n9867 & n22390;
  assign n25662 = n10434 & n22387;
  assign n25663 = ~n25661 & ~n25662;
  assign n25664 = ~n25660 & n25663;
  assign n25665 = n9870 & n22806;
  assign n25666 = n25664 & ~n25665;
  assign n25667 =  a[5]  & ~n25666;
  assign n25668 = ~n25666 & ~n25667;
  assign n25669 =  a[5]  & ~n25667;
  assign n25670 = ~n25668 & ~n25669;
  assign n25671 = n25010 & ~n25012;
  assign n25672 = ~n25013 & ~n25671;
  assign n25673 = ~n25670 & n25672;
  assign n25674 = ~n25670 & ~n25673;
  assign n25675 = n25672 & ~n25673;
  assign n25676 = ~n25674 & ~n25675;
  assign n25677 = ~n24997 & ~n25009;
  assign n25678 = ~n25008 & ~n25009;
  assign n25679 = ~n25677 & ~n25678;
  assign n25680 = n71 & n22387;
  assign n25681 = n9867 & n22393;
  assign n25682 = n10434 & n22390;
  assign n25683 = ~n25681 & ~n25682;
  assign n25684 = ~n25680 & n25683;
  assign n25685 = ~n9870 & n25684;
  assign n25686 = ~n22582 & n25684;
  assign n25687 = ~n25685 & ~n25686;
  assign n25688 =  a[5]  & ~n25687;
  assign n25689 = ~ a[5]  & n25687;
  assign n25690 = ~n25688 & ~n25689;
  assign n25691 = ~n25679 & ~n25690;
  assign n25692 = n71 & n22390;
  assign n25693 = n9867 & n22396;
  assign n25694 = n10434 & n22393;
  assign n25695 = ~n25693 & ~n25694;
  assign n25696 = ~n25692 & n25695;
  assign n25697 = n9870 & n22649;
  assign n25698 = n25696 & ~n25697;
  assign n25699 =  a[5]  & ~n25698;
  assign n25700 = ~n25698 & ~n25699;
  assign n25701 =  a[5]  & ~n25699;
  assign n25702 = ~n25700 & ~n25701;
  assign n25703 = ~n24981 & n24992;
  assign n25704 = ~n24993 & ~n25703;
  assign n25705 = ~n25702 & n25704;
  assign n25706 = ~n25702 & ~n25705;
  assign n25707 = n25704 & ~n25705;
  assign n25708 = ~n25706 & ~n25707;
  assign n25709 = n24978 & ~n24980;
  assign n25710 = ~n24981 & ~n25709;
  assign n25711 = n71 & n22393;
  assign n25712 = n9867 & n22399;
  assign n25713 = n10434 & n22396;
  assign n25714 = ~n25712 & ~n25713;
  assign n25715 = ~n25711 & n25714;
  assign n25716 = ~n9870 & n25715;
  assign n25717 = ~n22671 & n25715;
  assign n25718 = ~n25716 & ~n25717;
  assign n25719 =  a[5]  & ~n25718;
  assign n25720 = ~ a[5]  & n25718;
  assign n25721 = ~n25719 & ~n25720;
  assign n25722 = n25710 & ~n25721;
  assign n25723 = n10434 & ~n22406;
  assign n25724 = n71 & n22402;
  assign n25725 = ~n25723 & ~n25724;
  assign n25726 = n9870 & ~n22609;
  assign n25727 = n25725 & ~n25726;
  assign n25728 =  a[5]  & ~n25727;
  assign n25729 =  a[5]  & ~n25728;
  assign n25730 = ~n25727 & ~n25728;
  assign n25731 = ~n25729 & ~n25730;
  assign n25732 = ~n70 & ~n22406;
  assign n25733 =  a[5]  & ~n25732;
  assign n25734 = ~n25731 & n25733;
  assign n25735 = n71 & n22399;
  assign n25736 = n9867 & ~n22406;
  assign n25737 = n10434 & n22402;
  assign n25738 = ~n25736 & ~n25737;
  assign n25739 = ~n25735 & n25738;
  assign n25740 = ~n9870 & n25739;
  assign n25741 = n22625 & n25739;
  assign n25742 = ~n25740 & ~n25741;
  assign n25743 =  a[5]  & ~n25742;
  assign n25744 = ~ a[5]  & n25742;
  assign n25745 = ~n25743 & ~n25744;
  assign n25746 = n25734 & ~n25745;
  assign n25747 = n24979 & n25746;
  assign n25748 = n25746 & ~n25747;
  assign n25749 = n24979 & ~n25747;
  assign n25750 = ~n25748 & ~n25749;
  assign n25751 = n71 & n22396;
  assign n25752 = n9867 & n22402;
  assign n25753 = n10434 & n22399;
  assign n25754 = ~n25752 & ~n25753;
  assign n25755 = ~n25751 & n25754;
  assign n25756 = n9870 & n22595;
  assign n25757 = n25755 & ~n25756;
  assign n25758 =  a[5]  & ~n25757;
  assign n25759 =  a[5]  & ~n25758;
  assign n25760 = ~n25757 & ~n25758;
  assign n25761 = ~n25759 & ~n25760;
  assign n25762 = ~n25750 & ~n25761;
  assign n25763 = ~n25747 & ~n25762;
  assign n25764 = ~n25710 & n25721;
  assign n25765 = ~n25722 & ~n25764;
  assign n25766 = ~n25763 & n25765;
  assign n25767 = ~n25722 & ~n25766;
  assign n25768 = ~n25708 & ~n25767;
  assign n25769 = ~n25705 & ~n25768;
  assign n25770 = n25679 & n25690;
  assign n25771 = ~n25691 & ~n25770;
  assign n25772 = ~n25769 & n25771;
  assign n25773 = ~n25691 & ~n25772;
  assign n25774 = ~n25676 & ~n25773;
  assign n25775 = ~n25673 & ~n25774;
  assign n25776 = n25647 & ~n25659;
  assign n25777 = ~n25658 & ~n25659;
  assign n25778 = ~n25776 & ~n25777;
  assign n25779 = ~n25775 & ~n25778;
  assign n25780 = ~n25659 & ~n25779;
  assign n25781 = n25633 & ~n25645;
  assign n25782 = ~n25644 & ~n25645;
  assign n25783 = ~n25781 & ~n25782;
  assign n25784 = ~n25780 & ~n25783;
  assign n25785 = ~n25645 & ~n25784;
  assign n25786 = ~n25619 & n25630;
  assign n25787 = ~n25631 & ~n25786;
  assign n25788 = ~n25785 & n25787;
  assign n25789 = ~n25631 & ~n25788;
  assign n25790 = ~n25617 & ~n25789;
  assign n25791 = ~n25614 & ~n25790;
  assign n25792 = ~n25599 & ~n25791;
  assign n25793 = ~n25596 & ~n25792;
  assign n25794 = ~n25581 & ~n25793;
  assign n25795 = ~n25578 & ~n25794;
  assign n25796 = n25552 & ~n25564;
  assign n25797 = ~n25563 & ~n25564;
  assign n25798 = ~n25796 & ~n25797;
  assign n25799 = ~n25795 & ~n25798;
  assign n25800 = ~n25564 & ~n25799;
  assign n25801 = n25538 & ~n25550;
  assign n25802 = ~n25549 & ~n25550;
  assign n25803 = ~n25801 & ~n25802;
  assign n25804 = ~n25800 & ~n25803;
  assign n25805 = ~n25550 & ~n25804;
  assign n25806 = ~n25524 & n25535;
  assign n25807 = ~n25536 & ~n25806;
  assign n25808 = ~n25805 & n25807;
  assign n25809 = ~n25536 & ~n25808;
  assign n25810 = ~n25522 & ~n25809;
  assign n25811 = ~n25519 & ~n25810;
  assign n25812 = ~n25504 & ~n25811;
  assign n25813 = ~n25501 & ~n25812;
  assign n25814 = ~n25486 & ~n25813;
  assign n25815 = ~n25483 & ~n25814;
  assign n25816 = n25457 & ~n25469;
  assign n25817 = ~n25468 & ~n25469;
  assign n25818 = ~n25816 & ~n25817;
  assign n25819 = ~n25815 & ~n25818;
  assign n25820 = ~n25469 & ~n25819;
  assign n25821 = n25443 & ~n25455;
  assign n25822 = ~n25454 & ~n25455;
  assign n25823 = ~n25821 & ~n25822;
  assign n25824 = ~n25820 & ~n25823;
  assign n25825 = ~n25455 & ~n25824;
  assign n25826 = ~n25429 & n25440;
  assign n25827 = ~n25441 & ~n25826;
  assign n25828 = ~n25825 & n25827;
  assign n25829 = ~n25441 & ~n25828;
  assign n25830 = ~n25427 & ~n25829;
  assign n25831 = ~n25424 & ~n25830;
  assign n25832 = ~n25409 & ~n25831;
  assign n25833 = ~n25406 & ~n25832;
  assign n25834 = ~n25391 & ~n25833;
  assign n25835 = ~n25388 & ~n25834;
  assign n25836 = n25362 & ~n25374;
  assign n25837 = ~n25373 & ~n25374;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = ~n25835 & ~n25838;
  assign n25840 = ~n25374 & ~n25839;
  assign n25841 = ~n25348 & n25359;
  assign n25842 = ~n25360 & ~n25841;
  assign n25843 = ~n25840 & n25842;
  assign n25844 = ~n25360 & ~n25843;
  assign n25845 = ~n25346 & ~n25844;
  assign n25846 = ~n25343 & ~n25845;
  assign n25847 = ~n25328 & ~n25846;
  assign n25848 = ~n25325 & ~n25847;
  assign n25849 = ~n25307 & ~n25848;
  assign n25850 = ~n25304 & ~n25849;
  assign n25851 = n25287 & n25850;
  assign n25852 = ~n25287 & ~n25850;
  assign n25853 = ~n25851 & ~n25852;
  assign n25854 = ~n22284 & ~n22297;
  assign n25855 = ~n22275 & ~n22278;
  assign n25856 = ~n22270 & ~n22272;
  assign n25857 = n774 & n6716;
  assign n25858 = n1824 & n25857;
  assign n25859 = n3886 & n25858;
  assign n25860 = ~n619 & n25859;
  assign n25861 = ~n452 & n25860;
  assign n25862 = ~n1203 & n25861;
  assign n25863 = ~n237 & n25862;
  assign n25864 = n792 & n13063;
  assign n25865 = n3432 & n25864;
  assign n25866 = n3764 & n25865;
  assign n25867 = n3405 & n25866;
  assign n25868 = n1601 & n25867;
  assign n25869 = n25863 & n25868;
  assign n25870 = n2276 & n25869;
  assign n25871 = n1367 & n25870;
  assign n25872 = ~n364 & n25871;
  assign n25873 = ~n495 & n25872;
  assign n25874 = ~n296 & n25873;
  assign n25875 = ~n25856 & n25874;
  assign n25876 = n25856 & ~n25874;
  assign n25877 = ~n25875 & ~n25876;
  assign n25878 = n3020 & n13515;
  assign n25879 = n3028 & n13521;
  assign n25880 = n3023 & n13518;
  assign n25881 = n75 & n13541;
  assign n25882 = ~n25880 & ~n25881;
  assign n25883 = ~n25879 & n25882;
  assign n25884 = ~n25878 & n25883;
  assign n25885 = n25877 & ~n25884;
  assign n25886 = ~n25877 & n25884;
  assign n25887 = ~n25885 & ~n25886;
  assign n25888 = ~n25855 & n25887;
  assign n25889 = n25855 & ~n25887;
  assign n25890 = ~n25888 & ~n25889;
  assign n25891 = n3457 & n13633;
  assign n25892 = n3542 & n13597;
  assign n25893 = n3606 & n13630;
  assign n25894 = ~n25892 & ~n25893;
  assign n25895 = ~n25891 & n25894;
  assign n25896 = ~n3368 & n25895;
  assign n25897 = ~n13929 & n25895;
  assign n25898 = ~n25896 & ~n25897;
  assign n25899 =  a[29]  & ~n25898;
  assign n25900 = ~ a[29]  & n25898;
  assign n25901 = ~n25899 & ~n25900;
  assign n25902 = n25890 & ~n25901;
  assign n25903 = ~n25890 & n25901;
  assign n25904 = ~n25902 & ~n25903;
  assign n25905 = ~n25854 & n25904;
  assign n25906 = n25854 & ~n25904;
  assign n25907 = ~n25905 & ~n25906;
  assign n25908 = n3884 & ~n13438;
  assign n25909 = n3967 & ~n13627;
  assign n25910 = n4046 & n13941;
  assign n25911 = ~n25909 & ~n25910;
  assign n25912 = ~n25908 & n25911;
  assign n25913 = n4050 & n14028;
  assign n25914 = n25912 & ~n25913;
  assign n25915 =  a[26]  & ~n25914;
  assign n25916 =  a[26]  & ~n25915;
  assign n25917 = ~n25914 & ~n25915;
  assign n25918 = ~n25916 & ~n25917;
  assign n25919 = n25907 & ~n25918;
  assign n25920 = ~n25905 & ~n25919;
  assign n25921 = n75 & ~n13612;
  assign n25922 = n3020 & n13597;
  assign n25923 = n3023 & n13521;
  assign n25924 = n3028 & n13515;
  assign n25925 = ~n25923 & ~n25924;
  assign n25926 = ~n25922 & n25925;
  assign n25927 = ~n25921 & n25926;
  assign n25928 = n473 & n1047;
  assign n25929 = n3978 & n25928;
  assign n25930 = n3782 & n25929;
  assign n25931 = n13063 & n25930;
  assign n25932 = n1731 & n25931;
  assign n25933 = n2170 & n25932;
  assign n25934 = n3757 & n25933;
  assign n25935 = ~n746 & n25934;
  assign n25936 = ~n296 & n25935;
  assign n25937 = ~n173 & n25936;
  assign n25938 = ~n601 & n25937;
  assign n25939 = ~n245 & n25938;
  assign n25940 = ~n142 & n25939;
  assign n25941 = ~n25874 & n25940;
  assign n25942 = n25874 & ~n25940;
  assign n25943 = ~n25927 & ~n25942;
  assign n25944 = ~n25941 & n25943;
  assign n25945 = ~n25927 & ~n25944;
  assign n25946 = ~n25942 & ~n25944;
  assign n25947 = ~n25941 & n25946;
  assign n25948 = ~n25945 & ~n25947;
  assign n25949 = ~n25875 & ~n25885;
  assign n25950 = n25948 & n25949;
  assign n25951 = ~n25948 & ~n25949;
  assign n25952 = ~n25950 & ~n25951;
  assign n25953 = ~n25888 & ~n25902;
  assign n25954 = ~n25952 & n25953;
  assign n25955 = n25952 & ~n25953;
  assign n25956 = ~n25954 & ~n25955;
  assign n25957 = ~n3884 & ~n4046;
  assign n25958 = ~n13438 & ~n25957;
  assign n25959 = n3967 & n13941;
  assign n25960 = ~n25958 & ~n25959;
  assign n25961 = n4050 & ~n13951;
  assign n25962 = n25960 & ~n25961;
  assign n25963 =  a[26]  & ~n25962;
  assign n25964 = ~n25962 & ~n25963;
  assign n25965 =  a[26]  & ~n25963;
  assign n25966 = ~n25964 & ~n25965;
  assign n25967 = n3457 & ~n13627;
  assign n25968 = n3542 & n13630;
  assign n25969 = n3606 & n13633;
  assign n25970 = ~n25968 & ~n25969;
  assign n25971 = ~n25967 & n25970;
  assign n25972 = n3368 & ~n13654;
  assign n25973 = n25971 & ~n25972;
  assign n25974 =  a[29]  & ~n25973;
  assign n25975 =  a[29]  & ~n25974;
  assign n25976 = ~n25973 & ~n25974;
  assign n25977 = ~n25975 & ~n25976;
  assign n25978 = ~n25966 & ~n25977;
  assign n25979 = ~n25966 & ~n25978;
  assign n25980 = ~n25977 & ~n25978;
  assign n25981 = ~n25979 & ~n25980;
  assign n25982 = ~n25956 & n25981;
  assign n25983 = n25956 & ~n25981;
  assign n25984 = ~n25982 & ~n25983;
  assign n25985 = ~n25920 & n25984;
  assign n25986 = n25907 & ~n25919;
  assign n25987 = ~n25918 & ~n25919;
  assign n25988 = ~n25986 & ~n25987;
  assign n25989 = ~n22239 & ~n22300;
  assign n25990 = ~n22236 & ~n25989;
  assign n25991 = ~n25988 & ~n25990;
  assign n25992 = ~n25988 & ~n25991;
  assign n25993 = ~n25990 & ~n25991;
  assign n25994 = ~n25992 & ~n25993;
  assign n25995 = ~n22304 & ~n22307;
  assign n25996 = ~n25994 & ~n25995;
  assign n25997 = ~n25991 & ~n25996;
  assign n25998 = n25920 & ~n25984;
  assign n25999 = ~n25985 & ~n25998;
  assign n26000 = ~n25997 & n25999;
  assign n26001 = ~n25985 & ~n26000;
  assign n26002 = n75 & n13976;
  assign n26003 = n3020 & n13630;
  assign n26004 = n3023 & n13515;
  assign n26005 = n3028 & n13597;
  assign n26006 = ~n26004 & ~n26005;
  assign n26007 = ~n26003 & n26006;
  assign n26008 = ~n26002 & n26007;
  assign n26009 = ~n3967 & n25957;
  assign n26010 = ~n4050 & n26009;
  assign n26011 = ~n13438 & ~n26010;
  assign n26012 =  a[26]  & ~n26011;
  assign n26013 = ~ a[26]  & n26011;
  assign n26014 = ~n26012 & ~n26013;
  assign n26015 = n3873 & n3972;
  assign n26016 = ~n296 & n26015;
  assign n26017 = n4017 & n4040;
  assign n26018 = n2740 & n26017;
  assign n26019 = n26016 & n26018;
  assign n26020 = ~n328 & n26019;
  assign n26021 = ~n601 & n26020;
  assign n26022 = n25874 & n26021;
  assign n26023 = ~n25874 & ~n26021;
  assign n26024 = ~n26022 & ~n26023;
  assign n26025 = n26014 & n26024;
  assign n26026 = ~n26014 & ~n26024;
  assign n26027 = ~n26025 & ~n26026;
  assign n26028 = ~n25946 & n26027;
  assign n26029 = n25946 & ~n26027;
  assign n26030 = ~n26028 & ~n26029;
  assign n26031 = ~n26008 & n26030;
  assign n26032 = n26030 & ~n26031;
  assign n26033 = ~n26008 & ~n26031;
  assign n26034 = ~n26032 & ~n26033;
  assign n26035 = n3457 & n13941;
  assign n26036 = n3542 & n13633;
  assign n26037 = n3606 & ~n13627;
  assign n26038 = ~n26036 & ~n26037;
  assign n26039 = ~n26035 & n26038;
  assign n26040 = n3368 & n14136;
  assign n26041 = n26039 & ~n26040;
  assign n26042 =  a[29]  & ~n26041;
  assign n26043 =  a[29]  & ~n26042;
  assign n26044 = ~n26041 & ~n26042;
  assign n26045 = ~n26043 & ~n26044;
  assign n26046 = ~n26034 & ~n26045;
  assign n26047 = ~n26034 & ~n26046;
  assign n26048 = ~n26045 & ~n26046;
  assign n26049 = ~n26047 & ~n26048;
  assign n26050 = ~n25951 & ~n25955;
  assign n26051 = n26049 & n26050;
  assign n26052 = ~n26049 & ~n26050;
  assign n26053 = ~n26051 & ~n26052;
  assign n26054 = ~n25978 & ~n25983;
  assign n26055 = n26053 & ~n26054;
  assign n26056 = ~n26053 & n26054;
  assign n26057 = ~n26055 & ~n26056;
  assign n26058 = n26001 & ~n26057;
  assign n26059 = ~n26001 & n26057;
  assign n26060 = ~n26058 & ~n26059;
  assign n26061 = n11727 & n26060;
  assign n26062 = n25994 & n25995;
  assign n26063 = ~n25996 & ~n26062;
  assign n26064 = n11055 & n26063;
  assign n26065 = n25997 & ~n25999;
  assign n26066 = ~n26000 & ~n26065;
  assign n26067 = n11715 & n26066;
  assign n26068 = ~n26064 & ~n26067;
  assign n26069 = ~n26061 & n26068;
  assign n26070 = ~n11057 & n26069;
  assign n26071 = n26063 & n26066;
  assign n26072 = n22309 & n26063;
  assign n26073 = ~n22309 & ~n26063;
  assign n26074 = ~n22527 & ~n26073;
  assign n26075 = ~n26072 & n26074;
  assign n26076 = ~n26072 & ~n26075;
  assign n26077 = ~n26063 & ~n26066;
  assign n26078 = ~n26076 & ~n26077;
  assign n26079 = ~n26071 & n26078;
  assign n26080 = ~n26071 & ~n26079;
  assign n26081 = n26060 & n26066;
  assign n26082 = ~n26060 & ~n26066;
  assign n26083 = ~n26080 & ~n26082;
  assign n26084 = ~n26081 & n26083;
  assign n26085 = ~n26080 & ~n26084;
  assign n26086 = ~n26081 & ~n26084;
  assign n26087 = ~n26082 & n26086;
  assign n26088 = ~n26085 & ~n26087;
  assign n26089 = n26069 & n26088;
  assign n26090 = ~n26070 & ~n26089;
  assign n26091 =  a[2]  & ~n26090;
  assign n26092 = ~ a[2]  & n26090;
  assign n26093 = ~n26091 & ~n26092;
  assign n26094 = n25853 & ~n26093;
  assign n26095 = n25840 & ~n25842;
  assign n26096 = ~n25843 & ~n26095;
  assign n26097 = n25825 & ~n25827;
  assign n26098 = ~n25828 & ~n26097;
  assign n26099 = n25805 & ~n25807;
  assign n26100 = ~n25808 & ~n26099;
  assign n26101 = n25785 & ~n25787;
  assign n26102 = ~n25788 & ~n26101;
  assign n26103 = n25763 & ~n25765;
  assign n26104 = ~n25766 & ~n26103;
  assign n26105 = ~n25734 & n25745;
  assign n26106 = ~n25746 & ~n26105;
  assign n26107 = ~n11794 & ~n22406;
  assign n26108 = n11796 & ~n22625;
  assign n26109 = n11727 & n22399;
  assign n26110 = n11055 & ~n22406;
  assign n26111 = n11715 & n22402;
  assign n26112 = ~n26110 & ~n26111;
  assign n26113 = ~n26109 & n26112;
  assign n26114 =  a[2]  & ~n26113;
  assign n26115 = n11796 & ~n22609;
  assign n26116 = n11805 & ~n22406;
  assign n26117 = n11807 & n22402;
  assign n26118 =  a[2]  & ~n26117;
  assign n26119 = ~n26116 & n26118;
  assign n26120 = ~n26115 & n26119;
  assign n26121 = ~n26114 & n26120;
  assign n26122 = ~n26108 & n26121;
  assign n26123 = ~n26107 & n26122;
  assign n26124 = n25732 & n26123;
  assign n26125 = ~n25732 & ~n26123;
  assign n26126 = n11727 & n22396;
  assign n26127 = n11055 & n22402;
  assign n26128 = n11715 & n22399;
  assign n26129 = ~n26127 & ~n26128;
  assign n26130 = ~n26126 & n26129;
  assign n26131 = n11057 & n22595;
  assign n26132 = n26130 & ~n26131;
  assign n26133 = ~ a[2]  & ~n26132;
  assign n26134 =  a[2]  & n26132;
  assign n26135 = ~n26133 & ~n26134;
  assign n26136 = ~n26125 & ~n26135;
  assign n26137 = ~n26124 & ~n26136;
  assign n26138 = n11727 & n22393;
  assign n26139 = n11055 & n22399;
  assign n26140 = n11715 & n22396;
  assign n26141 = ~n26139 & ~n26140;
  assign n26142 = ~n26138 & n26141;
  assign n26143 = ~n11057 & n26142;
  assign n26144 = ~n22671 & n26142;
  assign n26145 = ~n26143 & ~n26144;
  assign n26146 =  a[2]  & ~n26145;
  assign n26147 = ~ a[2]  & n26145;
  assign n26148 = ~n26146 & ~n26147;
  assign n26149 = n26137 & n26148;
  assign n26150 = n25731 & ~n25733;
  assign n26151 = ~n25734 & ~n26150;
  assign n26152 = ~n26149 & n26151;
  assign n26153 = ~n26137 & ~n26148;
  assign n26154 = ~n26152 & ~n26153;
  assign n26155 = n26106 & ~n26154;
  assign n26156 = ~n26106 & n26154;
  assign n26157 = n11727 & n22390;
  assign n26158 = n11055 & n22396;
  assign n26159 = n11715 & n22393;
  assign n26160 = ~n26158 & ~n26159;
  assign n26161 = ~n26157 & n26160;
  assign n26162 = n11057 & n22649;
  assign n26163 = n26161 & ~n26162;
  assign n26164 = ~ a[2]  & ~n26163;
  assign n26165 =  a[2]  & n26163;
  assign n26166 = ~n26164 & ~n26165;
  assign n26167 = ~n26156 & ~n26166;
  assign n26168 = ~n26155 & ~n26167;
  assign n26169 = n11727 & n22387;
  assign n26170 = n11055 & n22393;
  assign n26171 = n11715 & n22390;
  assign n26172 = ~n26170 & ~n26171;
  assign n26173 = ~n26169 & n26172;
  assign n26174 = ~n11057 & n26173;
  assign n26175 = ~n22582 & n26173;
  assign n26176 = ~n26174 & ~n26175;
  assign n26177 =  a[2]  & ~n26176;
  assign n26178 = ~ a[2]  & n26176;
  assign n26179 = ~n26177 & ~n26178;
  assign n26180 = ~n26168 & ~n26179;
  assign n26181 = n26168 & n26179;
  assign n26182 = n25750 & n25761;
  assign n26183 = ~n25762 & ~n26182;
  assign n26184 = ~n26181 & n26183;
  assign n26185 = ~n26180 & ~n26184;
  assign n26186 = n26104 & ~n26185;
  assign n26187 = ~n26104 & n26185;
  assign n26188 = n11727 & n22384;
  assign n26189 = n11055 & n22390;
  assign n26190 = n11715 & n22387;
  assign n26191 = ~n26189 & ~n26190;
  assign n26192 = ~n26188 & n26191;
  assign n26193 = n11057 & n22806;
  assign n26194 = n26192 & ~n26193;
  assign n26195 = ~ a[2]  & ~n26194;
  assign n26196 =  a[2]  & n26194;
  assign n26197 = ~n26195 & ~n26196;
  assign n26198 = ~n26187 & ~n26197;
  assign n26199 = ~n26186 & ~n26198;
  assign n26200 = n11727 & n22380;
  assign n26201 = n11055 & n22387;
  assign n26202 = n11715 & n22384;
  assign n26203 = ~n26201 & ~n26202;
  assign n26204 = ~n26200 & n26203;
  assign n26205 = ~n11057 & n26204;
  assign n26206 = ~n22850 & n26204;
  assign n26207 = ~n26205 & ~n26206;
  assign n26208 =  a[2]  & ~n26207;
  assign n26209 = ~ a[2]  & n26207;
  assign n26210 = ~n26208 & ~n26209;
  assign n26211 = n26199 & n26210;
  assign n26212 = n25708 & n25767;
  assign n26213 = ~n25768 & ~n26212;
  assign n26214 = ~n26211 & n26213;
  assign n26215 = ~n26199 & ~n26210;
  assign n26216 = ~n26214 & ~n26215;
  assign n26217 = n11727 & n22377;
  assign n26218 = n11055 & n22384;
  assign n26219 = n11715 & n22380;
  assign n26220 = ~n26218 & ~n26219;
  assign n26221 = ~n26217 & n26220;
  assign n26222 = ~n11057 & n26221;
  assign n26223 = n22834 & n26221;
  assign n26224 = ~n26222 & ~n26223;
  assign n26225 =  a[2]  & ~n26224;
  assign n26226 = ~ a[2]  & n26224;
  assign n26227 = ~n26225 & ~n26226;
  assign n26228 = n26216 & n26227;
  assign n26229 = n25769 & ~n25771;
  assign n26230 = ~n25772 & ~n26229;
  assign n26231 = ~n26228 & n26230;
  assign n26232 = ~n26216 & ~n26227;
  assign n26233 = ~n26231 & ~n26232;
  assign n26234 = n11727 & n22374;
  assign n26235 = n11055 & n22380;
  assign n26236 = n11715 & n22377;
  assign n26237 = ~n26235 & ~n26236;
  assign n26238 = ~n26234 & n26237;
  assign n26239 = ~n11057 & n26238;
  assign n26240 = ~n22569 & n26238;
  assign n26241 = ~n26239 & ~n26240;
  assign n26242 =  a[2]  & ~n26241;
  assign n26243 = ~ a[2]  & n26241;
  assign n26244 = ~n26242 & ~n26243;
  assign n26245 = n26233 & n26244;
  assign n26246 = n25676 & n25773;
  assign n26247 = ~n25774 & ~n26246;
  assign n26248 = ~n26245 & n26247;
  assign n26249 = ~n26233 & ~n26244;
  assign n26250 = ~n26248 & ~n26249;
  assign n26251 = n25775 & ~n25777;
  assign n26252 = ~n25776 & n26251;
  assign n26253 = ~n25779 & ~n26252;
  assign n26254 = ~n26250 & n26253;
  assign n26255 = n26250 & ~n26253;
  assign n26256 = n11727 & n22371;
  assign n26257 = n11055 & n22377;
  assign n26258 = n11715 & n22374;
  assign n26259 = ~n26257 & ~n26258;
  assign n26260 = ~n26256 & n26259;
  assign n26261 = n11057 & n23025;
  assign n26262 = n26260 & ~n26261;
  assign n26263 = ~ a[2]  & ~n26262;
  assign n26264 =  a[2]  & n26262;
  assign n26265 = ~n26263 & ~n26264;
  assign n26266 = ~n26255 & ~n26265;
  assign n26267 = ~n26254 & ~n26266;
  assign n26268 = n25780 & ~n25782;
  assign n26269 = ~n25781 & n26268;
  assign n26270 = ~n25784 & ~n26269;
  assign n26271 = ~n26267 & n26270;
  assign n26272 = n26267 & ~n26270;
  assign n26273 = n11727 & n22368;
  assign n26274 = n11055 & n22374;
  assign n26275 = n11715 & n22371;
  assign n26276 = ~n26274 & ~n26275;
  assign n26277 = ~n26273 & n26276;
  assign n26278 = n11057 & n23006;
  assign n26279 = n26277 & ~n26278;
  assign n26280 = ~ a[2]  & ~n26279;
  assign n26281 =  a[2]  & n26279;
  assign n26282 = ~n26280 & ~n26281;
  assign n26283 = ~n26272 & ~n26282;
  assign n26284 = ~n26271 & ~n26283;
  assign n26285 = n26102 & ~n26284;
  assign n26286 = ~n26102 & n26284;
  assign n26287 = n11727 & n22365;
  assign n26288 = n11055 & n22371;
  assign n26289 = n11715 & n22368;
  assign n26290 = ~n26288 & ~n26289;
  assign n26291 = ~n26287 & n26290;
  assign n26292 = n11057 & ~n22993;
  assign n26293 = n26291 & ~n26292;
  assign n26294 = ~ a[2]  & ~n26293;
  assign n26295 =  a[2]  & n26293;
  assign n26296 = ~n26294 & ~n26295;
  assign n26297 = ~n26286 & ~n26296;
  assign n26298 = ~n26285 & ~n26297;
  assign n26299 = n11727 & n22362;
  assign n26300 = n11055 & n22368;
  assign n26301 = n11715 & n22365;
  assign n26302 = ~n26300 & ~n26301;
  assign n26303 = ~n26299 & n26302;
  assign n26304 = ~n11057 & n26303;
  assign n26305 = n23320 & n26303;
  assign n26306 = ~n26304 & ~n26305;
  assign n26307 =  a[2]  & ~n26306;
  assign n26308 = ~ a[2]  & n26306;
  assign n26309 = ~n26307 & ~n26308;
  assign n26310 = n26298 & n26309;
  assign n26311 = n25617 & n25789;
  assign n26312 = ~n25790 & ~n26311;
  assign n26313 = ~n26310 & n26312;
  assign n26314 = ~n26298 & ~n26309;
  assign n26315 = ~n26313 & ~n26314;
  assign n26316 = n11727 & n22359;
  assign n26317 = n11055 & n22365;
  assign n26318 = n11715 & n22362;
  assign n26319 = ~n26317 & ~n26318;
  assign n26320 = ~n26316 & n26319;
  assign n26321 = ~n11057 & n26320;
  assign n26322 = ~n23368 & n26320;
  assign n26323 = ~n26321 & ~n26322;
  assign n26324 =  a[2]  & ~n26323;
  assign n26325 = ~ a[2]  & n26323;
  assign n26326 = ~n26324 & ~n26325;
  assign n26327 = n26315 & n26326;
  assign n26328 = n25599 & n25791;
  assign n26329 = ~n25792 & ~n26328;
  assign n26330 = ~n26327 & n26329;
  assign n26331 = ~n26315 & ~n26326;
  assign n26332 = ~n26330 & ~n26331;
  assign n26333 = n11727 & n22356;
  assign n26334 = n11055 & n22362;
  assign n26335 = n11715 & n22359;
  assign n26336 = ~n26334 & ~n26335;
  assign n26337 = ~n26333 & n26336;
  assign n26338 = ~n11057 & n26337;
  assign n26339 = n23345 & n26337;
  assign n26340 = ~n26338 & ~n26339;
  assign n26341 =  a[2]  & ~n26340;
  assign n26342 = ~ a[2]  & n26340;
  assign n26343 = ~n26341 & ~n26342;
  assign n26344 = n26332 & n26343;
  assign n26345 = n25581 & n25793;
  assign n26346 = ~n25794 & ~n26345;
  assign n26347 = ~n26344 & n26346;
  assign n26348 = ~n26332 & ~n26343;
  assign n26349 = ~n26347 & ~n26348;
  assign n26350 = n25795 & ~n25797;
  assign n26351 = ~n25796 & n26350;
  assign n26352 = ~n25799 & ~n26351;
  assign n26353 = ~n26349 & n26352;
  assign n26354 = n26349 & ~n26352;
  assign n26355 = n11727 & n22353;
  assign n26356 = n11055 & n22359;
  assign n26357 = n11715 & n22356;
  assign n26358 = ~n26356 & ~n26357;
  assign n26359 = ~n26355 & n26358;
  assign n26360 = n11057 & ~n22556;
  assign n26361 = n26359 & ~n26360;
  assign n26362 = ~ a[2]  & ~n26361;
  assign n26363 =  a[2]  & n26361;
  assign n26364 = ~n26362 & ~n26363;
  assign n26365 = ~n26354 & ~n26364;
  assign n26366 = ~n26353 & ~n26365;
  assign n26367 = n25800 & ~n25802;
  assign n26368 = ~n25801 & n26367;
  assign n26369 = ~n25804 & ~n26368;
  assign n26370 = ~n26366 & n26369;
  assign n26371 = n26366 & ~n26369;
  assign n26372 = n11727 & n22350;
  assign n26373 = n11055 & n22356;
  assign n26374 = n11715 & n22353;
  assign n26375 = ~n26373 & ~n26374;
  assign n26376 = ~n26372 & n26375;
  assign n26377 = n11057 & n23672;
  assign n26378 = n26376 & ~n26377;
  assign n26379 = ~ a[2]  & ~n26378;
  assign n26380 =  a[2]  & n26378;
  assign n26381 = ~n26379 & ~n26380;
  assign n26382 = ~n26371 & ~n26381;
  assign n26383 = ~n26370 & ~n26382;
  assign n26384 = n26100 & ~n26383;
  assign n26385 = ~n26100 & n26383;
  assign n26386 = n11727 & n22347;
  assign n26387 = n11055 & n22353;
  assign n26388 = n11715 & n22350;
  assign n26389 = ~n26387 & ~n26388;
  assign n26390 = ~n26386 & n26389;
  assign n26391 = n11057 & ~n23659;
  assign n26392 = n26390 & ~n26391;
  assign n26393 = ~ a[2]  & ~n26392;
  assign n26394 =  a[2]  & n26392;
  assign n26395 = ~n26393 & ~n26394;
  assign n26396 = ~n26385 & ~n26395;
  assign n26397 = ~n26384 & ~n26396;
  assign n26398 = n11727 & n22344;
  assign n26399 = n11055 & n22350;
  assign n26400 = n11715 & n22347;
  assign n26401 = ~n26399 & ~n26400;
  assign n26402 = ~n26398 & n26401;
  assign n26403 = ~n11057 & n26402;
  assign n26404 = n23642 & n26402;
  assign n26405 = ~n26403 & ~n26404;
  assign n26406 =  a[2]  & ~n26405;
  assign n26407 = ~ a[2]  & n26405;
  assign n26408 = ~n26406 & ~n26407;
  assign n26409 = n26397 & n26408;
  assign n26410 = n25522 & n25809;
  assign n26411 = ~n25810 & ~n26410;
  assign n26412 = ~n26409 & n26411;
  assign n26413 = ~n26397 & ~n26408;
  assign n26414 = ~n26412 & ~n26413;
  assign n26415 = n11727 & n22341;
  assign n26416 = n11055 & n22347;
  assign n26417 = n11715 & n22344;
  assign n26418 = ~n26416 & ~n26417;
  assign n26419 = ~n26415 & n26418;
  assign n26420 = ~n11057 & n26419;
  assign n26421 = ~n24142 & n26419;
  assign n26422 = ~n26420 & ~n26421;
  assign n26423 =  a[2]  & ~n26422;
  assign n26424 = ~ a[2]  & n26422;
  assign n26425 = ~n26423 & ~n26424;
  assign n26426 = n26414 & n26425;
  assign n26427 = n25504 & n25811;
  assign n26428 = ~n25812 & ~n26427;
  assign n26429 = ~n26426 & n26428;
  assign n26430 = ~n26414 & ~n26425;
  assign n26431 = ~n26429 & ~n26430;
  assign n26432 = n11727 & n22338;
  assign n26433 = n11055 & n22344;
  assign n26434 = n11715 & n22341;
  assign n26435 = ~n26433 & ~n26434;
  assign n26436 = ~n26432 & n26435;
  assign n26437 = ~n11057 & n26436;
  assign n26438 = n24188 & n26436;
  assign n26439 = ~n26437 & ~n26438;
  assign n26440 =  a[2]  & ~n26439;
  assign n26441 = ~ a[2]  & n26439;
  assign n26442 = ~n26440 & ~n26441;
  assign n26443 = n26431 & n26442;
  assign n26444 = n25486 & n25813;
  assign n26445 = ~n25814 & ~n26444;
  assign n26446 = ~n26443 & n26445;
  assign n26447 = ~n26431 & ~n26442;
  assign n26448 = ~n26446 & ~n26447;
  assign n26449 = n25815 & ~n25817;
  assign n26450 = ~n25816 & n26449;
  assign n26451 = ~n25819 & ~n26450;
  assign n26452 = ~n26448 & n26451;
  assign n26453 = n26448 & ~n26451;
  assign n26454 = n11727 & n22335;
  assign n26455 = n11055 & n22341;
  assign n26456 = n11715 & n22338;
  assign n26457 = ~n26455 & ~n26456;
  assign n26458 = ~n26454 & n26457;
  assign n26459 = n11057 & ~n24167;
  assign n26460 = n26458 & ~n26459;
  assign n26461 = ~ a[2]  & ~n26460;
  assign n26462 =  a[2]  & n26460;
  assign n26463 = ~n26461 & ~n26462;
  assign n26464 = ~n26453 & ~n26463;
  assign n26465 = ~n26452 & ~n26464;
  assign n26466 = n25820 & ~n25822;
  assign n26467 = ~n25821 & n26466;
  assign n26468 = ~n25824 & ~n26467;
  assign n26469 = ~n26465 & n26468;
  assign n26470 = n26465 & ~n26468;
  assign n26471 = n11727 & n22332;
  assign n26472 = n11055 & n22338;
  assign n26473 = n11715 & n22335;
  assign n26474 = ~n26472 & ~n26473;
  assign n26475 = ~n26471 & n26474;
  assign n26476 = n11057 & n22542;
  assign n26477 = n26475 & ~n26476;
  assign n26478 = ~ a[2]  & ~n26477;
  assign n26479 =  a[2]  & n26477;
  assign n26480 = ~n26478 & ~n26479;
  assign n26481 = ~n26470 & ~n26480;
  assign n26482 = ~n26469 & ~n26481;
  assign n26483 = n26098 & ~n26482;
  assign n26484 = ~n26098 & n26482;
  assign n26485 = n11727 & n22329;
  assign n26486 = n11055 & n22335;
  assign n26487 = n11715 & n22332;
  assign n26488 = ~n26486 & ~n26487;
  assign n26489 = ~n26485 & n26488;
  assign n26490 = n11057 & ~n24633;
  assign n26491 = n26489 & ~n26490;
  assign n26492 = ~ a[2]  & ~n26491;
  assign n26493 =  a[2]  & n26491;
  assign n26494 = ~n26492 & ~n26493;
  assign n26495 = ~n26484 & ~n26494;
  assign n26496 = ~n26483 & ~n26495;
  assign n26497 = n11727 & n22326;
  assign n26498 = n11055 & n22332;
  assign n26499 = n11715 & n22329;
  assign n26500 = ~n26498 & ~n26499;
  assign n26501 = ~n26497 & n26500;
  assign n26502 = ~n11057 & n26501;
  assign n26503 = n24616 & n26501;
  assign n26504 = ~n26502 & ~n26503;
  assign n26505 =  a[2]  & ~n26504;
  assign n26506 = ~ a[2]  & n26504;
  assign n26507 = ~n26505 & ~n26506;
  assign n26508 = n26496 & n26507;
  assign n26509 = n25427 & n25829;
  assign n26510 = ~n25830 & ~n26509;
  assign n26511 = ~n26508 & n26510;
  assign n26512 = ~n26496 & ~n26507;
  assign n26513 = ~n26511 & ~n26512;
  assign n26514 = n11727 & n22323;
  assign n26515 = n11055 & n22329;
  assign n26516 = n11715 & n22326;
  assign n26517 = ~n26515 & ~n26516;
  assign n26518 = ~n26514 & n26517;
  assign n26519 = ~n11057 & n26518;
  assign n26520 = ~n24599 & n26518;
  assign n26521 = ~n26519 & ~n26520;
  assign n26522 =  a[2]  & ~n26521;
  assign n26523 = ~ a[2]  & n26521;
  assign n26524 = ~n26522 & ~n26523;
  assign n26525 = n26513 & n26524;
  assign n26526 = n25409 & n25831;
  assign n26527 = ~n25832 & ~n26526;
  assign n26528 = ~n26525 & n26527;
  assign n26529 = ~n26513 & ~n26524;
  assign n26530 = ~n26528 & ~n26529;
  assign n26531 = n11727 & n22320;
  assign n26532 = n11055 & n22326;
  assign n26533 = n11715 & n22323;
  assign n26534 = ~n26532 & ~n26533;
  assign n26535 = ~n26531 & n26534;
  assign n26536 = ~n11057 & n26535;
  assign n26537 = n25270 & n26535;
  assign n26538 = ~n26536 & ~n26537;
  assign n26539 =  a[2]  & ~n26538;
  assign n26540 = ~ a[2]  & n26538;
  assign n26541 = ~n26539 & ~n26540;
  assign n26542 = n26530 & n26541;
  assign n26543 = n25391 & n25833;
  assign n26544 = ~n25834 & ~n26543;
  assign n26545 = ~n26542 & n26544;
  assign n26546 = ~n26530 & ~n26541;
  assign n26547 = ~n26545 & ~n26546;
  assign n26548 = n25835 & ~n25837;
  assign n26549 = ~n25836 & n26548;
  assign n26550 = ~n25839 & ~n26549;
  assign n26551 = ~n26547 & n26550;
  assign n26552 = n26547 & ~n26550;
  assign n26553 = n11727 & n22312;
  assign n26554 = n11055 & n22323;
  assign n26555 = n11715 & n22320;
  assign n26556 = ~n26554 & ~n26555;
  assign n26557 = ~n26553 & n26556;
  assign n26558 = n11057 & ~n25315;
  assign n26559 = n26557 & ~n26558;
  assign n26560 = ~ a[2]  & ~n26559;
  assign n26561 =  a[2]  & n26559;
  assign n26562 = ~n26560 & ~n26561;
  assign n26563 = ~n26552 & ~n26562;
  assign n26564 = ~n26551 & ~n26563;
  assign n26565 = n26096 & ~n26564;
  assign n26566 = ~n26096 & n26564;
  assign n26567 = n11727 & n22315;
  assign n26568 = n11055 & n22320;
  assign n26569 = n11715 & n22312;
  assign n26570 = ~n26568 & ~n26569;
  assign n26571 = ~n26567 & n26570;
  assign n26572 = n11057 & n25294;
  assign n26573 = n26571 & ~n26572;
  assign n26574 = ~ a[2]  & ~n26573;
  assign n26575 =  a[2]  & n26573;
  assign n26576 = ~n26574 & ~n26575;
  assign n26577 = ~n26566 & ~n26576;
  assign n26578 = ~n26565 & ~n26577;
  assign n26579 = n11727 & n22309;
  assign n26580 = n11055 & n22312;
  assign n26581 = n11715 & n22315;
  assign n26582 = ~n26580 & ~n26581;
  assign n26583 = ~n26579 & n26582;
  assign n26584 = ~n11057 & n26583;
  assign n26585 = n22529 & n26583;
  assign n26586 = ~n26584 & ~n26585;
  assign n26587 =  a[2]  & ~n26586;
  assign n26588 = ~ a[2]  & n26586;
  assign n26589 = ~n26587 & ~n26588;
  assign n26590 = n26578 & n26589;
  assign n26591 = n25346 & n25844;
  assign n26592 = ~n25845 & ~n26591;
  assign n26593 = ~n26590 & n26592;
  assign n26594 = ~n26578 & ~n26589;
  assign n26595 = ~n26593 & ~n26594;
  assign n26596 = n11727 & n26063;
  assign n26597 = n11055 & n22315;
  assign n26598 = n11715 & n22309;
  assign n26599 = ~n26597 & ~n26598;
  assign n26600 = ~n26596 & n26599;
  assign n26601 = ~n11057 & n26600;
  assign n26602 = ~n22527 & ~n26075;
  assign n26603 = ~n26073 & n26076;
  assign n26604 = ~n26602 & ~n26603;
  assign n26605 = n26600 & n26604;
  assign n26606 = ~n26601 & ~n26605;
  assign n26607 =  a[2]  & ~n26606;
  assign n26608 = ~ a[2]  & n26606;
  assign n26609 = ~n26607 & ~n26608;
  assign n26610 = n26595 & n26609;
  assign n26611 = n25328 & n25846;
  assign n26612 = ~n25847 & ~n26611;
  assign n26613 = ~n26610 & n26612;
  assign n26614 = ~n26595 & ~n26609;
  assign n26615 = ~n26613 & ~n26614;
  assign n26616 = n11727 & n26066;
  assign n26617 = n11055 & n22309;
  assign n26618 = n11715 & n26063;
  assign n26619 = ~n26617 & ~n26618;
  assign n26620 = ~n26616 & n26619;
  assign n26621 = ~n11057 & n26620;
  assign n26622 = ~n26076 & ~n26079;
  assign n26623 = ~n26077 & n26080;
  assign n26624 = ~n26622 & ~n26623;
  assign n26625 = n26620 & n26624;
  assign n26626 = ~n26621 & ~n26625;
  assign n26627 =  a[2]  & ~n26626;
  assign n26628 = ~ a[2]  & n26626;
  assign n26629 = ~n26627 & ~n26628;
  assign n26630 = n26615 & n26629;
  assign n26631 = n25307 & n25848;
  assign n26632 = ~n25849 & ~n26631;
  assign n26633 = ~n26630 & n26632;
  assign n26634 = ~n26615 & ~n26629;
  assign n26635 = ~n26633 & ~n26634;
  assign n26636 = n25853 & ~n26094;
  assign n26637 = ~n26093 & ~n26094;
  assign n26638 = ~n26636 & ~n26637;
  assign n26639 = ~n26635 & ~n26638;
  assign n26640 = ~n26094 & ~n26639;
  assign n26641 = n71 & n26063;
  assign n26642 = n9867 & n22315;
  assign n26643 = n10434 & n22309;
  assign n26644 = ~n26642 & ~n26643;
  assign n26645 = ~n26641 & n26644;
  assign n26646 = n9870 & ~n26604;
  assign n26647 = n26645 & ~n26646;
  assign n26648 =  a[5]  & ~n26647;
  assign n26649 = ~n26647 & ~n26648;
  assign n26650 =  a[5]  & ~n26648;
  assign n26651 = ~n26649 & ~n26650;
  assign n26652 = ~n25276 & ~n25280;
  assign n26653 = n7983 & n22326;
  assign n26654 = n7291 & n22332;
  assign n26655 = n7632 & n22329;
  assign n26656 = ~n26654 & ~n26655;
  assign n26657 = ~n26653 & n26656;
  assign n26658 = n7294 & ~n24616;
  assign n26659 = n26657 & ~n26658;
  assign n26660 =  a[11]  & ~n26659;
  assign n26661 = ~n26659 & ~n26660;
  assign n26662 =  a[11]  & ~n26660;
  assign n26663 = ~n26661 & ~n26662;
  assign n26664 = ~n25246 & ~n25250;
  assign n26665 = n6233 & n22344;
  assign n26666 = n5663 & n22350;
  assign n26667 = n5939 & n22347;
  assign n26668 = ~n26666 & ~n26667;
  assign n26669 = ~n26665 & n26668;
  assign n26670 = n5666 & ~n23642;
  assign n26671 = n26669 & ~n26670;
  assign n26672 =  a[17]  & ~n26671;
  assign n26673 = ~n26671 & ~n26672;
  assign n26674 =  a[17]  & ~n26672;
  assign n26675 = ~n26673 & ~n26674;
  assign n26676 = ~n25219 & ~n25223;
  assign n26677 = n4694 & n22362;
  assign n26678 = n4533 & n22368;
  assign n26679 = n4604 & n22365;
  assign n26680 = ~n26678 & ~n26679;
  assign n26681 = ~n26677 & n26680;
  assign n26682 = n4536 & ~n23320;
  assign n26683 = n26681 & ~n26682;
  assign n26684 =  a[23]  & ~n26683;
  assign n26685 = ~n26683 & ~n26684;
  assign n26686 =  a[23]  & ~n26684;
  assign n26687 = ~n26685 & ~n26686;
  assign n26688 = ~n25192 & ~n25196;
  assign n26689 = n3457 & n22380;
  assign n26690 = n3542 & n22387;
  assign n26691 = n3606 & n22384;
  assign n26692 = ~n26690 & ~n26691;
  assign n26693 = ~n26689 & n26692;
  assign n26694 = n3368 & n22850;
  assign n26695 = n26693 & ~n26694;
  assign n26696 =  a[29]  & ~n26695;
  assign n26697 = ~n26695 & ~n26696;
  assign n26698 =  a[29]  & ~n26696;
  assign n26699 = ~n26697 & ~n26698;
  assign n26700 = ~n25165 & ~n25169;
  assign n26701 = n12397 & n13789;
  assign n26702 = n4771 & n26701;
  assign n26703 = n1887 & n26702;
  assign n26704 = n790 & n26703;
  assign n26705 = n13677 & n26704;
  assign n26706 = n4311 & n26705;
  assign n26707 = n3155 & n26706;
  assign n26708 = n244 & n26707;
  assign n26709 = n933 & n26708;
  assign n26710 = n1237 & n26709;
  assign n26711 = n116 & n26710;
  assign n26712 = ~n1101 & n26711;
  assign n26713 = ~n422 & n26712;
  assign n26714 = ~n493 & n26713;
  assign n26715 = ~n428 & n26714;
  assign n26716 = n3020 & n22390;
  assign n26717 = n3028 & n22393;
  assign n26718 = n3023 & n22396;
  assign n26719 = n75 & n22649;
  assign n26720 = ~n26718 & ~n26719;
  assign n26721 = ~n26717 & n26720;
  assign n26722 = ~n26716 & n26721;
  assign n26723 = ~n26715 & ~n26722;
  assign n26724 = ~n26715 & ~n26723;
  assign n26725 = ~n26722 & ~n26723;
  assign n26726 = ~n26724 & ~n26725;
  assign n26727 = ~n26700 & ~n26726;
  assign n26728 = ~n26700 & ~n26727;
  assign n26729 = ~n26726 & ~n26727;
  assign n26730 = ~n26728 & ~n26729;
  assign n26731 = ~n26699 & ~n26730;
  assign n26732 = ~n26699 & ~n26731;
  assign n26733 = ~n26730 & ~n26731;
  assign n26734 = ~n26732 & ~n26733;
  assign n26735 = ~n25173 & ~n25179;
  assign n26736 = n26734 & n26735;
  assign n26737 = ~n26734 & ~n26735;
  assign n26738 = ~n26736 & ~n26737;
  assign n26739 = n3884 & n22371;
  assign n26740 = n3967 & n22377;
  assign n26741 = n4046 & n22374;
  assign n26742 = ~n26740 & ~n26741;
  assign n26743 = ~n26739 & n26742;
  assign n26744 = ~n4050 & n26743;
  assign n26745 = ~n23025 & n26743;
  assign n26746 = ~n26744 & ~n26745;
  assign n26747 =  a[26]  & ~n26746;
  assign n26748 = ~ a[26]  & n26746;
  assign n26749 = ~n26747 & ~n26748;
  assign n26750 = n26738 & ~n26749;
  assign n26751 = n26738 & ~n26750;
  assign n26752 = ~n26749 & ~n26750;
  assign n26753 = ~n26751 & ~n26752;
  assign n26754 = ~n26688 & ~n26753;
  assign n26755 = ~n26688 & ~n26754;
  assign n26756 = ~n26753 & ~n26754;
  assign n26757 = ~n26755 & ~n26756;
  assign n26758 = ~n26687 & ~n26757;
  assign n26759 = ~n26687 & ~n26758;
  assign n26760 = ~n26757 & ~n26758;
  assign n26761 = ~n26759 & ~n26760;
  assign n26762 = ~n25200 & ~n25206;
  assign n26763 = n26761 & n26762;
  assign n26764 = ~n26761 & ~n26762;
  assign n26765 = ~n26763 & ~n26764;
  assign n26766 = n5496 & n22353;
  assign n26767 = n4935 & n22359;
  assign n26768 = n5407 & n22356;
  assign n26769 = ~n26767 & ~n26768;
  assign n26770 = ~n26766 & n26769;
  assign n26771 = ~n4938 & n26770;
  assign n26772 = n22556 & n26770;
  assign n26773 = ~n26771 & ~n26772;
  assign n26774 =  a[20]  & ~n26773;
  assign n26775 = ~ a[20]  & n26773;
  assign n26776 = ~n26774 & ~n26775;
  assign n26777 = n26765 & ~n26776;
  assign n26778 = n26765 & ~n26777;
  assign n26779 = ~n26776 & ~n26777;
  assign n26780 = ~n26778 & ~n26779;
  assign n26781 = ~n26676 & ~n26780;
  assign n26782 = ~n26676 & ~n26781;
  assign n26783 = ~n26780 & ~n26781;
  assign n26784 = ~n26782 & ~n26783;
  assign n26785 = ~n26675 & ~n26784;
  assign n26786 = ~n26675 & ~n26785;
  assign n26787 = ~n26784 & ~n26785;
  assign n26788 = ~n26786 & ~n26787;
  assign n26789 = ~n25227 & ~n25233;
  assign n26790 = n26788 & n26789;
  assign n26791 = ~n26788 & ~n26789;
  assign n26792 = ~n26790 & ~n26791;
  assign n26793 = n7101 & n22335;
  assign n26794 = n6402 & n22341;
  assign n26795 = n6951 & n22338;
  assign n26796 = ~n26794 & ~n26795;
  assign n26797 = ~n26793 & n26796;
  assign n26798 = ~n6397 & n26797;
  assign n26799 = n24167 & n26797;
  assign n26800 = ~n26798 & ~n26799;
  assign n26801 =  a[14]  & ~n26800;
  assign n26802 = ~ a[14]  & n26800;
  assign n26803 = ~n26801 & ~n26802;
  assign n26804 = n26792 & ~n26803;
  assign n26805 = n26792 & ~n26804;
  assign n26806 = ~n26803 & ~n26804;
  assign n26807 = ~n26805 & ~n26806;
  assign n26808 = ~n26664 & ~n26807;
  assign n26809 = ~n26664 & ~n26808;
  assign n26810 = ~n26807 & ~n26808;
  assign n26811 = ~n26809 & ~n26810;
  assign n26812 = ~n26663 & ~n26811;
  assign n26813 = ~n26663 & ~n26812;
  assign n26814 = ~n26811 & ~n26812;
  assign n26815 = ~n26813 & ~n26814;
  assign n26816 = ~n25254 & ~n25260;
  assign n26817 = n26815 & n26816;
  assign n26818 = ~n26815 & ~n26816;
  assign n26819 = ~n26817 & ~n26818;
  assign n26820 = n9331 & n22312;
  assign n26821 = n8418 & n22323;
  assign n26822 = n8860 & n22320;
  assign n26823 = ~n26821 & ~n26822;
  assign n26824 = ~n26820 & n26823;
  assign n26825 = ~n8421 & n26824;
  assign n26826 = n25315 & n26824;
  assign n26827 = ~n26825 & ~n26826;
  assign n26828 =  a[8]  & ~n26827;
  assign n26829 = ~ a[8]  & n26827;
  assign n26830 = ~n26828 & ~n26829;
  assign n26831 = n26819 & ~n26830;
  assign n26832 = n26819 & ~n26831;
  assign n26833 = ~n26830 & ~n26831;
  assign n26834 = ~n26832 & ~n26833;
  assign n26835 = ~n26652 & ~n26834;
  assign n26836 = ~n26652 & ~n26835;
  assign n26837 = ~n26834 & ~n26835;
  assign n26838 = ~n26836 & ~n26837;
  assign n26839 = ~n26651 & ~n26838;
  assign n26840 = ~n26651 & ~n26839;
  assign n26841 = ~n26838 & ~n26839;
  assign n26842 = ~n26840 & ~n26841;
  assign n26843 = ~n25284 & ~n25852;
  assign n26844 = n26842 & n26843;
  assign n26845 = ~n26842 & ~n26843;
  assign n26846 = ~n26844 & ~n26845;
  assign n26847 = ~n26055 & ~n26059;
  assign n26848 = ~n26046 & ~n26052;
  assign n26849 = n75 & n13929;
  assign n26850 = n3020 & n13633;
  assign n26851 = n3023 & n13597;
  assign n26852 = n3028 & n13630;
  assign n26853 = ~n26851 & ~n26852;
  assign n26854 = ~n26850 & n26853;
  assign n26855 = ~n26849 & n26854;
  assign n26856 = ~n26023 & ~n26025;
  assign n26857 = n4030 & n4511;
  assign n26858 = n26016 & n26857;
  assign n26859 = ~n328 & n26858;
  assign n26860 = ~n26856 & n26859;
  assign n26861 = n26856 & ~n26859;
  assign n26862 = ~n26860 & ~n26861;
  assign n26863 = ~n26855 & n26862;
  assign n26864 = ~n26855 & ~n26863;
  assign n26865 = n26862 & ~n26863;
  assign n26866 = ~n26864 & ~n26865;
  assign n26867 = ~n26028 & ~n26031;
  assign n26868 = n26866 & n26867;
  assign n26869 = ~n26866 & ~n26867;
  assign n26870 = ~n26868 & ~n26869;
  assign n26871 = n3457 & ~n13438;
  assign n26872 = n3542 & ~n13627;
  assign n26873 = n3606 & n13941;
  assign n26874 = ~n26872 & ~n26873;
  assign n26875 = ~n26871 & n26874;
  assign n26876 = ~n3368 & n26875;
  assign n26877 = ~n14028 & n26875;
  assign n26878 = ~n26876 & ~n26877;
  assign n26879 =  a[29]  & ~n26878;
  assign n26880 = ~ a[29]  & n26878;
  assign n26881 = ~n26879 & ~n26880;
  assign n26882 = n26870 & ~n26881;
  assign n26883 = ~n26870 & n26881;
  assign n26884 = ~n26882 & ~n26883;
  assign n26885 = ~n26848 & n26884;
  assign n26886 = n26848 & ~n26884;
  assign n26887 = ~n26885 & ~n26886;
  assign n26888 = ~n26847 & n26887;
  assign n26889 = n26847 & ~n26887;
  assign n26890 = ~n26888 & ~n26889;
  assign n26891 = n11727 & n26890;
  assign n26892 = n11055 & n26066;
  assign n26893 = n11715 & n26060;
  assign n26894 = ~n26892 & ~n26893;
  assign n26895 = ~n26891 & n26894;
  assign n26896 = ~n11057 & n26895;
  assign n26897 = n26060 & n26890;
  assign n26898 = ~n26060 & ~n26890;
  assign n26899 = ~n26086 & ~n26898;
  assign n26900 = ~n26897 & n26899;
  assign n26901 = ~n26086 & ~n26900;
  assign n26902 = ~n26897 & ~n26900;
  assign n26903 = ~n26898 & n26902;
  assign n26904 = ~n26901 & ~n26903;
  assign n26905 = n26895 & n26904;
  assign n26906 = ~n26896 & ~n26905;
  assign n26907 =  a[2]  & ~n26906;
  assign n26908 = ~ a[2]  & n26906;
  assign n26909 = ~n26907 & ~n26908;
  assign n26910 = n26846 & ~n26909;
  assign n26911 = ~n26846 & n26909;
  assign n26912 = ~n26910 & ~n26911;
  assign n26913 = ~n26640 & n26912;
  assign n26914 = n26640 & ~n26912;
  assign n26915 = ~n26913 & ~n26914;
  assign n26916 = ~n26635 & ~n26639;
  assign n26917 = ~n26638 & ~n26639;
  assign n26918 = ~n26916 & ~n26917;
  assign n26919 = n26915 & n26918;
  assign n26920 = ~n26915 & ~n26918;
  assign  result[0]  = n26919 | n26920;
  assign n26922 = n26915 & ~n26918;
  assign n26923 = ~n26910 & ~n26913;
  assign n26924 = n71 & n26066;
  assign n26925 = n9867 & n22309;
  assign n26926 = n10434 & n26063;
  assign n26927 = ~n26925 & ~n26926;
  assign n26928 = ~n26924 & n26927;
  assign n26929 = n9870 & ~n26624;
  assign n26930 = n26928 & ~n26929;
  assign n26931 =  a[5]  & ~n26930;
  assign n26932 = ~n26930 & ~n26931;
  assign n26933 =  a[5]  & ~n26931;
  assign n26934 = ~n26932 & ~n26933;
  assign n26935 = ~n26831 & ~n26835;
  assign n26936 = n7983 & n22323;
  assign n26937 = n7291 & n22329;
  assign n26938 = n7632 & n22326;
  assign n26939 = ~n26937 & ~n26938;
  assign n26940 = ~n26936 & n26939;
  assign n26941 = n7294 & n24599;
  assign n26942 = n26940 & ~n26941;
  assign n26943 =  a[11]  & ~n26942;
  assign n26944 = ~n26942 & ~n26943;
  assign n26945 =  a[11]  & ~n26943;
  assign n26946 = ~n26944 & ~n26945;
  assign n26947 = ~n26804 & ~n26808;
  assign n26948 = n6233 & n22341;
  assign n26949 = n5663 & n22347;
  assign n26950 = n5939 & n22344;
  assign n26951 = ~n26949 & ~n26950;
  assign n26952 = ~n26948 & n26951;
  assign n26953 = n5666 & n24142;
  assign n26954 = n26952 & ~n26953;
  assign n26955 =  a[17]  & ~n26954;
  assign n26956 = ~n26954 & ~n26955;
  assign n26957 =  a[17]  & ~n26955;
  assign n26958 = ~n26956 & ~n26957;
  assign n26959 = ~n26777 & ~n26781;
  assign n26960 = n4694 & n22359;
  assign n26961 = n4533 & n22365;
  assign n26962 = n4604 & n22362;
  assign n26963 = ~n26961 & ~n26962;
  assign n26964 = ~n26960 & n26963;
  assign n26965 = n4536 & n23368;
  assign n26966 = n26964 & ~n26965;
  assign n26967 =  a[23]  & ~n26966;
  assign n26968 = ~n26966 & ~n26967;
  assign n26969 =  a[23]  & ~n26967;
  assign n26970 = ~n26968 & ~n26969;
  assign n26971 = ~n26750 & ~n26754;
  assign n26972 = ~n26731 & ~n26737;
  assign n26973 = ~n26723 & ~n26727;
  assign n26974 = n1603 & n3514;
  assign n26975 = n2025 & n26974;
  assign n26976 = n6628 & n26975;
  assign n26977 = n14544 & n26976;
  assign n26978 = n6755 & n26977;
  assign n26979 = n2979 & n26978;
  assign n26980 = n3544 & n26979;
  assign n26981 = n1575 & n26980;
  assign n26982 = n2583 & n26981;
  assign n26983 = n1237 & n26982;
  assign n26984 = n2405 & n26983;
  assign n26985 = n1522 & n26984;
  assign n26986 = ~n1246 & n26985;
  assign n26987 = ~n330 & n26986;
  assign n26988 = ~n296 & n26987;
  assign n26989 = ~n372 & n26988;
  assign n26990 = ~n932 & n26989;
  assign n26991 = ~n771 & n26990;
  assign n26992 = n3020 & n22387;
  assign n26993 = n3028 & n22390;
  assign n26994 = n3023 & n22393;
  assign n26995 = n75 & n22582;
  assign n26996 = ~n26994 & ~n26995;
  assign n26997 = ~n26993 & n26996;
  assign n26998 = ~n26992 & n26997;
  assign n26999 = ~n26991 & ~n26998;
  assign n27000 = ~n26991 & ~n26999;
  assign n27001 = ~n26998 & ~n26999;
  assign n27002 = ~n27000 & ~n27001;
  assign n27003 = ~n26973 & ~n27002;
  assign n27004 = ~n26973 & ~n27003;
  assign n27005 = ~n27002 & ~n27003;
  assign n27006 = ~n27004 & ~n27005;
  assign n27007 = n3457 & n22377;
  assign n27008 = n3542 & n22384;
  assign n27009 = n3606 & n22380;
  assign n27010 = ~n27008 & ~n27009;
  assign n27011 = ~n27007 & n27010;
  assign n27012 = ~n3368 & n27011;
  assign n27013 = n22834 & n27011;
  assign n27014 = ~n27012 & ~n27013;
  assign n27015 =  a[29]  & ~n27014;
  assign n27016 = ~ a[29]  & n27014;
  assign n27017 = ~n27015 & ~n27016;
  assign n27018 = ~n27006 & ~n27017;
  assign n27019 = n27006 & n27017;
  assign n27020 = ~n27018 & ~n27019;
  assign n27021 = ~n26972 & n27020;
  assign n27022 = n26972 & ~n27020;
  assign n27023 = ~n27021 & ~n27022;
  assign n27024 = n3884 & n22368;
  assign n27025 = n3967 & n22374;
  assign n27026 = n4046 & n22371;
  assign n27027 = ~n27025 & ~n27026;
  assign n27028 = ~n27024 & n27027;
  assign n27029 = ~n4050 & n27028;
  assign n27030 = ~n23006 & n27028;
  assign n27031 = ~n27029 & ~n27030;
  assign n27032 =  a[26]  & ~n27031;
  assign n27033 = ~ a[26]  & n27031;
  assign n27034 = ~n27032 & ~n27033;
  assign n27035 = n27023 & ~n27034;
  assign n27036 = n27023 & ~n27035;
  assign n27037 = ~n27034 & ~n27035;
  assign n27038 = ~n27036 & ~n27037;
  assign n27039 = ~n26971 & ~n27038;
  assign n27040 = ~n26971 & ~n27039;
  assign n27041 = ~n27038 & ~n27039;
  assign n27042 = ~n27040 & ~n27041;
  assign n27043 = ~n26970 & ~n27042;
  assign n27044 = ~n26970 & ~n27043;
  assign n27045 = ~n27042 & ~n27043;
  assign n27046 = ~n27044 & ~n27045;
  assign n27047 = ~n26758 & ~n26764;
  assign n27048 = n27046 & n27047;
  assign n27049 = ~n27046 & ~n27047;
  assign n27050 = ~n27048 & ~n27049;
  assign n27051 = n5496 & n22350;
  assign n27052 = n4935 & n22356;
  assign n27053 = n5407 & n22353;
  assign n27054 = ~n27052 & ~n27053;
  assign n27055 = ~n27051 & n27054;
  assign n27056 = ~n4938 & n27055;
  assign n27057 = ~n23672 & n27055;
  assign n27058 = ~n27056 & ~n27057;
  assign n27059 =  a[20]  & ~n27058;
  assign n27060 = ~ a[20]  & n27058;
  assign n27061 = ~n27059 & ~n27060;
  assign n27062 = n27050 & ~n27061;
  assign n27063 = n27050 & ~n27062;
  assign n27064 = ~n27061 & ~n27062;
  assign n27065 = ~n27063 & ~n27064;
  assign n27066 = ~n26959 & ~n27065;
  assign n27067 = ~n26959 & ~n27066;
  assign n27068 = ~n27065 & ~n27066;
  assign n27069 = ~n27067 & ~n27068;
  assign n27070 = ~n26958 & ~n27069;
  assign n27071 = ~n26958 & ~n27070;
  assign n27072 = ~n27069 & ~n27070;
  assign n27073 = ~n27071 & ~n27072;
  assign n27074 = ~n26785 & ~n26791;
  assign n27075 = n27073 & n27074;
  assign n27076 = ~n27073 & ~n27074;
  assign n27077 = ~n27075 & ~n27076;
  assign n27078 = n7101 & n22332;
  assign n27079 = n6402 & n22338;
  assign n27080 = n6951 & n22335;
  assign n27081 = ~n27079 & ~n27080;
  assign n27082 = ~n27078 & n27081;
  assign n27083 = ~n6397 & n27082;
  assign n27084 = ~n22542 & n27082;
  assign n27085 = ~n27083 & ~n27084;
  assign n27086 =  a[14]  & ~n27085;
  assign n27087 = ~ a[14]  & n27085;
  assign n27088 = ~n27086 & ~n27087;
  assign n27089 = n27077 & ~n27088;
  assign n27090 = n27077 & ~n27089;
  assign n27091 = ~n27088 & ~n27089;
  assign n27092 = ~n27090 & ~n27091;
  assign n27093 = ~n26947 & ~n27092;
  assign n27094 = ~n26947 & ~n27093;
  assign n27095 = ~n27092 & ~n27093;
  assign n27096 = ~n27094 & ~n27095;
  assign n27097 = ~n26946 & ~n27096;
  assign n27098 = ~n26946 & ~n27097;
  assign n27099 = ~n27096 & ~n27097;
  assign n27100 = ~n27098 & ~n27099;
  assign n27101 = ~n26812 & ~n26818;
  assign n27102 = n27100 & n27101;
  assign n27103 = ~n27100 & ~n27101;
  assign n27104 = ~n27102 & ~n27103;
  assign n27105 = n9331 & n22315;
  assign n27106 = n8418 & n22320;
  assign n27107 = n8860 & n22312;
  assign n27108 = ~n27106 & ~n27107;
  assign n27109 = ~n27105 & n27108;
  assign n27110 = ~n8421 & n27109;
  assign n27111 = ~n25294 & n27109;
  assign n27112 = ~n27110 & ~n27111;
  assign n27113 =  a[8]  & ~n27112;
  assign n27114 = ~ a[8]  & n27112;
  assign n27115 = ~n27113 & ~n27114;
  assign n27116 = n27104 & ~n27115;
  assign n27117 = n27104 & ~n27116;
  assign n27118 = ~n27115 & ~n27116;
  assign n27119 = ~n27117 & ~n27118;
  assign n27120 = ~n26935 & ~n27119;
  assign n27121 = ~n26935 & ~n27120;
  assign n27122 = ~n27119 & ~n27120;
  assign n27123 = ~n27121 & ~n27122;
  assign n27124 = ~n26934 & ~n27123;
  assign n27125 = ~n26934 & ~n27124;
  assign n27126 = ~n27123 & ~n27124;
  assign n27127 = ~n27125 & ~n27126;
  assign n27128 = ~n26839 & ~n26845;
  assign n27129 = n27127 & n27128;
  assign n27130 = ~n27127 & ~n27128;
  assign n27131 = ~n27129 & ~n27130;
  assign n27132 = ~n26885 & ~n26888;
  assign n27133 = ~n26869 & ~n26882;
  assign n27134 = ~n26860 & ~n26863;
  assign n27135 = n3856 & n4514;
  assign n27136 = n26859 & ~n27135;
  assign n27137 = ~n26859 & n27135;
  assign n27138 = ~n27134 & ~n27137;
  assign n27139 = ~n27136 & n27138;
  assign n27140 = ~n27134 & ~n27139;
  assign n27141 = ~n27137 & ~n27139;
  assign n27142 = ~n27136 & n27141;
  assign n27143 = ~n27140 & ~n27142;
  assign n27144 = ~n3457 & ~n3606;
  assign n27145 = ~n13438 & ~n27144;
  assign n27146 = n3542 & n13941;
  assign n27147 = ~n27145 & ~n27146;
  assign n27148 = n3368 & ~n13951;
  assign n27149 = n27147 & ~n27148;
  assign n27150 =  a[29]  & ~n27149;
  assign n27151 = ~n27149 & ~n27150;
  assign n27152 =  a[29]  & ~n27150;
  assign n27153 = ~n27151 & ~n27152;
  assign n27154 = n75 & ~n13654;
  assign n27155 = n3020 & ~n13627;
  assign n27156 = n3023 & n13630;
  assign n27157 = n3028 & n13633;
  assign n27158 = ~n27156 & ~n27157;
  assign n27159 = ~n27155 & n27158;
  assign n27160 = ~n27154 & n27159;
  assign n27161 = ~n27153 & ~n27160;
  assign n27162 = ~n27153 & ~n27161;
  assign n27163 = ~n27160 & ~n27161;
  assign n27164 = ~n27162 & ~n27163;
  assign n27165 = ~n27143 & n27164;
  assign n27166 = n27143 & ~n27164;
  assign n27167 = ~n27165 & ~n27166;
  assign n27168 = ~n27133 & ~n27167;
  assign n27169 = n27133 & n27167;
  assign n27170 = ~n27168 & ~n27169;
  assign n27171 = ~n27132 & n27170;
  assign n27172 = n27132 & ~n27170;
  assign n27173 = ~n27171 & ~n27172;
  assign n27174 = n11727 & n27173;
  assign n27175 = n11055 & n26060;
  assign n27176 = n11715 & n26890;
  assign n27177 = ~n27175 & ~n27176;
  assign n27178 = ~n27174 & n27177;
  assign n27179 = ~n11057 & n27178;
  assign n27180 = ~n26890 & ~n27173;
  assign n27181 = n26890 & n27173;
  assign n27182 = ~n27180 & ~n27181;
  assign n27183 = ~n26902 & n27182;
  assign n27184 = n26902 & ~n27182;
  assign n27185 = ~n27183 & ~n27184;
  assign n27186 = n27178 & ~n27185;
  assign n27187 = ~n27179 & ~n27186;
  assign n27188 =  a[2]  & ~n27187;
  assign n27189 = ~ a[2]  & n27187;
  assign n27190 = ~n27188 & ~n27189;
  assign n27191 = n27131 & ~n27190;
  assign n27192 = ~n27131 & n27190;
  assign n27193 = ~n27191 & ~n27192;
  assign n27194 = ~n26923 & n27193;
  assign n27195 = n26923 & ~n27193;
  assign n27196 = ~n27194 & ~n27195;
  assign n27197 = n26922 & n27196;
  assign n27198 = ~n26922 & ~n27196;
  assign  result[1]  = ~n27197 & ~n27198;
  assign n27200 = ~n27191 & ~n27194;
  assign n27201 = n71 & n26060;
  assign n27202 = n9867 & n26063;
  assign n27203 = n10434 & n26066;
  assign n27204 = ~n27202 & ~n27203;
  assign n27205 = ~n27201 & n27204;
  assign n27206 = n9870 & ~n26088;
  assign n27207 = n27205 & ~n27206;
  assign n27208 =  a[5]  & ~n27207;
  assign n27209 = ~n27207 & ~n27208;
  assign n27210 =  a[5]  & ~n27208;
  assign n27211 = ~n27209 & ~n27210;
  assign n27212 = ~n27116 & ~n27120;
  assign n27213 = n7983 & n22320;
  assign n27214 = n7291 & n22326;
  assign n27215 = n7632 & n22323;
  assign n27216 = ~n27214 & ~n27215;
  assign n27217 = ~n27213 & n27216;
  assign n27218 = n7294 & ~n25270;
  assign n27219 = n27217 & ~n27218;
  assign n27220 =  a[11]  & ~n27219;
  assign n27221 = ~n27219 & ~n27220;
  assign n27222 =  a[11]  & ~n27220;
  assign n27223 = ~n27221 & ~n27222;
  assign n27224 = ~n27089 & ~n27093;
  assign n27225 = n6233 & n22338;
  assign n27226 = n5663 & n22344;
  assign n27227 = n5939 & n22341;
  assign n27228 = ~n27226 & ~n27227;
  assign n27229 = ~n27225 & n27228;
  assign n27230 = n5666 & ~n24188;
  assign n27231 = n27229 & ~n27230;
  assign n27232 =  a[17]  & ~n27231;
  assign n27233 = ~n27231 & ~n27232;
  assign n27234 =  a[17]  & ~n27232;
  assign n27235 = ~n27233 & ~n27234;
  assign n27236 = ~n27062 & ~n27066;
  assign n27237 = n4694 & n22356;
  assign n27238 = n4533 & n22362;
  assign n27239 = n4604 & n22359;
  assign n27240 = ~n27238 & ~n27239;
  assign n27241 = ~n27237 & n27240;
  assign n27242 = n4536 & ~n23345;
  assign n27243 = n27241 & ~n27242;
  assign n27244 =  a[23]  & ~n27243;
  assign n27245 = ~n27243 & ~n27244;
  assign n27246 =  a[23]  & ~n27244;
  assign n27247 = ~n27245 & ~n27246;
  assign n27248 = ~n27035 & ~n27039;
  assign n27249 = ~n27018 & ~n27021;
  assign n27250 = ~n26999 & ~n27003;
  assign n27251 = n13827 & n14561;
  assign n27252 = n6717 & n27251;
  assign n27253 = n2410 & n27252;
  assign n27254 = n616 & n27253;
  assign n27255 = n3180 & n27254;
  assign n27256 = n3191 & n27255;
  assign n27257 = n1600 & n27256;
  assign n27258 = n1479 & n27257;
  assign n27259 = n1844 & n27258;
  assign n27260 = n515 & n27259;
  assign n27261 = n1726 & n27260;
  assign n27262 = n1269 & n27261;
  assign n27263 = ~n107 & n27262;
  assign n27264 = ~n490 & n27263;
  assign n27265 = ~n286 & n27264;
  assign n27266 = ~n245 & n27265;
  assign n27267 = ~n470 & n27266;
  assign n27268 = n3020 & n22384;
  assign n27269 = n3028 & n22387;
  assign n27270 = n3023 & n22390;
  assign n27271 = n75 & n22806;
  assign n27272 = ~n27270 & ~n27271;
  assign n27273 = ~n27269 & n27272;
  assign n27274 = ~n27268 & n27273;
  assign n27275 = ~n27267 & ~n27274;
  assign n27276 = ~n27267 & ~n27275;
  assign n27277 = ~n27274 & ~n27275;
  assign n27278 = ~n27276 & ~n27277;
  assign n27279 = ~n27250 & ~n27278;
  assign n27280 = ~n27250 & ~n27279;
  assign n27281 = ~n27278 & ~n27279;
  assign n27282 = ~n27280 & ~n27281;
  assign n27283 = n3457 & n22374;
  assign n27284 = n3542 & n22380;
  assign n27285 = n3606 & n22377;
  assign n27286 = ~n27284 & ~n27285;
  assign n27287 = ~n27283 & n27286;
  assign n27288 = ~n3368 & n27287;
  assign n27289 = ~n22569 & n27287;
  assign n27290 = ~n27288 & ~n27289;
  assign n27291 =  a[29]  & ~n27290;
  assign n27292 = ~ a[29]  & n27290;
  assign n27293 = ~n27291 & ~n27292;
  assign n27294 = ~n27282 & ~n27293;
  assign n27295 = n27282 & n27293;
  assign n27296 = ~n27294 & ~n27295;
  assign n27297 = ~n27249 & n27296;
  assign n27298 = n27249 & ~n27296;
  assign n27299 = ~n27297 & ~n27298;
  assign n27300 = n3884 & n22365;
  assign n27301 = n3967 & n22371;
  assign n27302 = n4046 & n22368;
  assign n27303 = ~n27301 & ~n27302;
  assign n27304 = ~n27300 & n27303;
  assign n27305 = ~n4050 & n27304;
  assign n27306 = n22993 & n27304;
  assign n27307 = ~n27305 & ~n27306;
  assign n27308 =  a[26]  & ~n27307;
  assign n27309 = ~ a[26]  & n27307;
  assign n27310 = ~n27308 & ~n27309;
  assign n27311 = n27299 & ~n27310;
  assign n27312 = n27299 & ~n27311;
  assign n27313 = ~n27310 & ~n27311;
  assign n27314 = ~n27312 & ~n27313;
  assign n27315 = ~n27248 & ~n27314;
  assign n27316 = ~n27248 & ~n27315;
  assign n27317 = ~n27314 & ~n27315;
  assign n27318 = ~n27316 & ~n27317;
  assign n27319 = ~n27247 & ~n27318;
  assign n27320 = ~n27247 & ~n27319;
  assign n27321 = ~n27318 & ~n27319;
  assign n27322 = ~n27320 & ~n27321;
  assign n27323 = ~n27043 & ~n27049;
  assign n27324 = n27322 & n27323;
  assign n27325 = ~n27322 & ~n27323;
  assign n27326 = ~n27324 & ~n27325;
  assign n27327 = n5496 & n22347;
  assign n27328 = n4935 & n22353;
  assign n27329 = n5407 & n22350;
  assign n27330 = ~n27328 & ~n27329;
  assign n27331 = ~n27327 & n27330;
  assign n27332 = ~n4938 & n27331;
  assign n27333 = n23659 & n27331;
  assign n27334 = ~n27332 & ~n27333;
  assign n27335 =  a[20]  & ~n27334;
  assign n27336 = ~ a[20]  & n27334;
  assign n27337 = ~n27335 & ~n27336;
  assign n27338 = n27326 & ~n27337;
  assign n27339 = n27326 & ~n27338;
  assign n27340 = ~n27337 & ~n27338;
  assign n27341 = ~n27339 & ~n27340;
  assign n27342 = ~n27236 & ~n27341;
  assign n27343 = ~n27236 & ~n27342;
  assign n27344 = ~n27341 & ~n27342;
  assign n27345 = ~n27343 & ~n27344;
  assign n27346 = ~n27235 & ~n27345;
  assign n27347 = ~n27235 & ~n27346;
  assign n27348 = ~n27345 & ~n27346;
  assign n27349 = ~n27347 & ~n27348;
  assign n27350 = ~n27070 & ~n27076;
  assign n27351 = n27349 & n27350;
  assign n27352 = ~n27349 & ~n27350;
  assign n27353 = ~n27351 & ~n27352;
  assign n27354 = n7101 & n22329;
  assign n27355 = n6402 & n22335;
  assign n27356 = n6951 & n22332;
  assign n27357 = ~n27355 & ~n27356;
  assign n27358 = ~n27354 & n27357;
  assign n27359 = ~n6397 & n27358;
  assign n27360 = n24633 & n27358;
  assign n27361 = ~n27359 & ~n27360;
  assign n27362 =  a[14]  & ~n27361;
  assign n27363 = ~ a[14]  & n27361;
  assign n27364 = ~n27362 & ~n27363;
  assign n27365 = n27353 & ~n27364;
  assign n27366 = n27353 & ~n27365;
  assign n27367 = ~n27364 & ~n27365;
  assign n27368 = ~n27366 & ~n27367;
  assign n27369 = ~n27224 & ~n27368;
  assign n27370 = ~n27224 & ~n27369;
  assign n27371 = ~n27368 & ~n27369;
  assign n27372 = ~n27370 & ~n27371;
  assign n27373 = ~n27223 & ~n27372;
  assign n27374 = ~n27223 & ~n27373;
  assign n27375 = ~n27372 & ~n27373;
  assign n27376 = ~n27374 & ~n27375;
  assign n27377 = ~n27097 & ~n27103;
  assign n27378 = n27376 & n27377;
  assign n27379 = ~n27376 & ~n27377;
  assign n27380 = ~n27378 & ~n27379;
  assign n27381 = n9331 & n22309;
  assign n27382 = n8418 & n22312;
  assign n27383 = n8860 & n22315;
  assign n27384 = ~n27382 & ~n27383;
  assign n27385 = ~n27381 & n27384;
  assign n27386 = ~n8421 & n27385;
  assign n27387 = n22529 & n27385;
  assign n27388 = ~n27386 & ~n27387;
  assign n27389 =  a[8]  & ~n27388;
  assign n27390 = ~ a[8]  & n27388;
  assign n27391 = ~n27389 & ~n27390;
  assign n27392 = n27380 & ~n27391;
  assign n27393 = n27380 & ~n27392;
  assign n27394 = ~n27391 & ~n27392;
  assign n27395 = ~n27393 & ~n27394;
  assign n27396 = ~n27212 & ~n27395;
  assign n27397 = ~n27212 & ~n27396;
  assign n27398 = ~n27395 & ~n27396;
  assign n27399 = ~n27397 & ~n27398;
  assign n27400 = ~n27211 & ~n27399;
  assign n27401 = ~n27211 & ~n27400;
  assign n27402 = ~n27399 & ~n27400;
  assign n27403 = ~n27401 & ~n27402;
  assign n27404 = ~n27124 & ~n27130;
  assign n27405 = n27403 & n27404;
  assign n27406 = ~n27403 & ~n27404;
  assign n27407 = ~n27405 & ~n27406;
  assign n27408 = ~n27168 & ~n27171;
  assign n27409 = ~n27143 & ~n27164;
  assign n27410 = ~n27161 & ~n27409;
  assign n27411 = n75 & n14136;
  assign n27412 = n3020 & n13941;
  assign n27413 = n3023 & n13633;
  assign n27414 = n3028 & ~n13627;
  assign n27415 = ~n27413 & ~n27414;
  assign n27416 = ~n27412 & n27415;
  assign n27417 = ~n27411 & n27416;
  assign n27418 = ~n3542 & ~n3606;
  assign n27419 = n3367 & n27418;
  assign n27420 = ~n13438 & ~n27419;
  assign n27421 =  a[29]  & ~n27420;
  assign n27422 = ~ a[29]  & n27420;
  assign n27423 = ~n27421 & ~n27422;
  assign n27424 = n13056 & n27135;
  assign n27425 = ~n13056 & ~n27135;
  assign n27426 = ~n27424 & ~n27425;
  assign n27427 = n27423 & n27426;
  assign n27428 = ~n27423 & ~n27426;
  assign n27429 = ~n27427 & ~n27428;
  assign n27430 = ~n27417 & n27429;
  assign n27431 = n27429 & ~n27430;
  assign n27432 = ~n27417 & ~n27430;
  assign n27433 = ~n27431 & ~n27432;
  assign n27434 = ~n27141 & ~n27433;
  assign n27435 = n27141 & n27433;
  assign n27436 = ~n27434 & ~n27435;
  assign n27437 = ~n27410 & n27436;
  assign n27438 = n27410 & ~n27436;
  assign n27439 = ~n27437 & ~n27438;
  assign n27440 = ~n27408 & n27439;
  assign n27441 = n27408 & ~n27439;
  assign n27442 = ~n27440 & ~n27441;
  assign n27443 = n11727 & n27442;
  assign n27444 = n11055 & n26890;
  assign n27445 = n11715 & n27173;
  assign n27446 = ~n27444 & ~n27445;
  assign n27447 = ~n27443 & n27446;
  assign n27448 = ~n11057 & n27447;
  assign n27449 = ~n27181 & ~n27183;
  assign n27450 = ~n27173 & ~n27442;
  assign n27451 = n27173 & n27442;
  assign n27452 = ~n27450 & ~n27451;
  assign n27453 = ~n27449 & n27452;
  assign n27454 = n27449 & ~n27452;
  assign n27455 = ~n27453 & ~n27454;
  assign n27456 = n27447 & ~n27455;
  assign n27457 = ~n27448 & ~n27456;
  assign n27458 =  a[2]  & ~n27457;
  assign n27459 = ~ a[2]  & n27457;
  assign n27460 = ~n27458 & ~n27459;
  assign n27461 = n27407 & ~n27460;
  assign n27462 = ~n27407 & n27460;
  assign n27463 = ~n27461 & ~n27462;
  assign n27464 = ~n27200 & n27463;
  assign n27465 = n27200 & ~n27463;
  assign n27466 = ~n27464 & ~n27465;
  assign n27467 = n27197 & n27466;
  assign n27468 = ~n27197 & ~n27466;
  assign  result[2]  = ~n27467 & ~n27468;
  assign n27470 = ~n27461 & ~n27464;
  assign n27471 = n71 & n26890;
  assign n27472 = n9867 & n26066;
  assign n27473 = n10434 & n26060;
  assign n27474 = ~n27472 & ~n27473;
  assign n27475 = ~n27471 & n27474;
  assign n27476 = n9870 & ~n26904;
  assign n27477 = n27475 & ~n27476;
  assign n27478 =  a[5]  & ~n27477;
  assign n27479 = ~n27477 & ~n27478;
  assign n27480 =  a[5]  & ~n27478;
  assign n27481 = ~n27479 & ~n27480;
  assign n27482 = ~n27392 & ~n27396;
  assign n27483 = n7983 & n22312;
  assign n27484 = n7291 & n22323;
  assign n27485 = n7632 & n22320;
  assign n27486 = ~n27484 & ~n27485;
  assign n27487 = ~n27483 & n27486;
  assign n27488 = n7294 & ~n25315;
  assign n27489 = n27487 & ~n27488;
  assign n27490 =  a[11]  & ~n27489;
  assign n27491 = ~n27489 & ~n27490;
  assign n27492 =  a[11]  & ~n27490;
  assign n27493 = ~n27491 & ~n27492;
  assign n27494 = ~n27365 & ~n27369;
  assign n27495 = n6233 & n22335;
  assign n27496 = n5663 & n22341;
  assign n27497 = n5939 & n22338;
  assign n27498 = ~n27496 & ~n27497;
  assign n27499 = ~n27495 & n27498;
  assign n27500 = n5666 & ~n24167;
  assign n27501 = n27499 & ~n27500;
  assign n27502 =  a[17]  & ~n27501;
  assign n27503 = ~n27501 & ~n27502;
  assign n27504 =  a[17]  & ~n27502;
  assign n27505 = ~n27503 & ~n27504;
  assign n27506 = ~n27338 & ~n27342;
  assign n27507 = n4694 & n22353;
  assign n27508 = n4533 & n22359;
  assign n27509 = n4604 & n22356;
  assign n27510 = ~n27508 & ~n27509;
  assign n27511 = ~n27507 & n27510;
  assign n27512 = n4536 & ~n22556;
  assign n27513 = n27511 & ~n27512;
  assign n27514 =  a[23]  & ~n27513;
  assign n27515 = ~n27513 & ~n27514;
  assign n27516 =  a[23]  & ~n27514;
  assign n27517 = ~n27515 & ~n27516;
  assign n27518 = ~n27311 & ~n27315;
  assign n27519 = ~n27294 & ~n27297;
  assign n27520 = ~n27275 & ~n27279;
  assign n27521 = n156 & n2466;
  assign n27522 = n2993 & n27521;
  assign n27523 = n1721 & n1737;
  assign n27524 = n27522 & n27523;
  assign n27525 = n2410 & n27524;
  assign n27526 = n4769 & n27525;
  assign n27527 = n15743 & n27526;
  assign n27528 = n6732 & n27527;
  assign n27529 = n6769 & n27528;
  assign n27530 = n2229 & n27529;
  assign n27531 = n510 & n27530;
  assign n27532 = n1826 & n27531;
  assign n27533 = n1182 & n27532;
  assign n27534 = ~n191 & n27533;
  assign n27535 = ~n340 & n27534;
  assign n27536 = n3020 & n22380;
  assign n27537 = n3028 & n22384;
  assign n27538 = n3023 & n22387;
  assign n27539 = n75 & n22850;
  assign n27540 = ~n27538 & ~n27539;
  assign n27541 = ~n27537 & n27540;
  assign n27542 = ~n27536 & n27541;
  assign n27543 = ~n27535 & ~n27542;
  assign n27544 = ~n27535 & ~n27543;
  assign n27545 = ~n27542 & ~n27543;
  assign n27546 = ~n27544 & ~n27545;
  assign n27547 = ~n27520 & ~n27546;
  assign n27548 = ~n27520 & ~n27547;
  assign n27549 = ~n27546 & ~n27547;
  assign n27550 = ~n27548 & ~n27549;
  assign n27551 = n3457 & n22371;
  assign n27552 = n3542 & n22377;
  assign n27553 = n3606 & n22374;
  assign n27554 = ~n27552 & ~n27553;
  assign n27555 = ~n27551 & n27554;
  assign n27556 = ~n3368 & n27555;
  assign n27557 = ~n23025 & n27555;
  assign n27558 = ~n27556 & ~n27557;
  assign n27559 =  a[29]  & ~n27558;
  assign n27560 = ~ a[29]  & n27558;
  assign n27561 = ~n27559 & ~n27560;
  assign n27562 = ~n27550 & ~n27561;
  assign n27563 = n27550 & n27561;
  assign n27564 = ~n27562 & ~n27563;
  assign n27565 = ~n27519 & n27564;
  assign n27566 = n27519 & ~n27564;
  assign n27567 = ~n27565 & ~n27566;
  assign n27568 = n3884 & n22362;
  assign n27569 = n3967 & n22368;
  assign n27570 = n4046 & n22365;
  assign n27571 = ~n27569 & ~n27570;
  assign n27572 = ~n27568 & n27571;
  assign n27573 = ~n4050 & n27572;
  assign n27574 = n23320 & n27572;
  assign n27575 = ~n27573 & ~n27574;
  assign n27576 =  a[26]  & ~n27575;
  assign n27577 = ~ a[26]  & n27575;
  assign n27578 = ~n27576 & ~n27577;
  assign n27579 = n27567 & ~n27578;
  assign n27580 = n27567 & ~n27579;
  assign n27581 = ~n27578 & ~n27579;
  assign n27582 = ~n27580 & ~n27581;
  assign n27583 = ~n27518 & ~n27582;
  assign n27584 = ~n27518 & ~n27583;
  assign n27585 = ~n27582 & ~n27583;
  assign n27586 = ~n27584 & ~n27585;
  assign n27587 = ~n27517 & ~n27586;
  assign n27588 = ~n27517 & ~n27587;
  assign n27589 = ~n27586 & ~n27587;
  assign n27590 = ~n27588 & ~n27589;
  assign n27591 = ~n27319 & ~n27325;
  assign n27592 = n27590 & n27591;
  assign n27593 = ~n27590 & ~n27591;
  assign n27594 = ~n27592 & ~n27593;
  assign n27595 = n5496 & n22344;
  assign n27596 = n4935 & n22350;
  assign n27597 = n5407 & n22347;
  assign n27598 = ~n27596 & ~n27597;
  assign n27599 = ~n27595 & n27598;
  assign n27600 = ~n4938 & n27599;
  assign n27601 = n23642 & n27599;
  assign n27602 = ~n27600 & ~n27601;
  assign n27603 =  a[20]  & ~n27602;
  assign n27604 = ~ a[20]  & n27602;
  assign n27605 = ~n27603 & ~n27604;
  assign n27606 = n27594 & ~n27605;
  assign n27607 = n27594 & ~n27606;
  assign n27608 = ~n27605 & ~n27606;
  assign n27609 = ~n27607 & ~n27608;
  assign n27610 = ~n27506 & ~n27609;
  assign n27611 = ~n27506 & ~n27610;
  assign n27612 = ~n27609 & ~n27610;
  assign n27613 = ~n27611 & ~n27612;
  assign n27614 = ~n27505 & ~n27613;
  assign n27615 = ~n27505 & ~n27614;
  assign n27616 = ~n27613 & ~n27614;
  assign n27617 = ~n27615 & ~n27616;
  assign n27618 = ~n27346 & ~n27352;
  assign n27619 = n27617 & n27618;
  assign n27620 = ~n27617 & ~n27618;
  assign n27621 = ~n27619 & ~n27620;
  assign n27622 = n7101 & n22326;
  assign n27623 = n6402 & n22332;
  assign n27624 = n6951 & n22329;
  assign n27625 = ~n27623 & ~n27624;
  assign n27626 = ~n27622 & n27625;
  assign n27627 = ~n6397 & n27626;
  assign n27628 = n24616 & n27626;
  assign n27629 = ~n27627 & ~n27628;
  assign n27630 =  a[14]  & ~n27629;
  assign n27631 = ~ a[14]  & n27629;
  assign n27632 = ~n27630 & ~n27631;
  assign n27633 = n27621 & ~n27632;
  assign n27634 = n27621 & ~n27633;
  assign n27635 = ~n27632 & ~n27633;
  assign n27636 = ~n27634 & ~n27635;
  assign n27637 = ~n27494 & ~n27636;
  assign n27638 = ~n27494 & ~n27637;
  assign n27639 = ~n27636 & ~n27637;
  assign n27640 = ~n27638 & ~n27639;
  assign n27641 = ~n27493 & ~n27640;
  assign n27642 = ~n27493 & ~n27641;
  assign n27643 = ~n27640 & ~n27641;
  assign n27644 = ~n27642 & ~n27643;
  assign n27645 = ~n27373 & ~n27379;
  assign n27646 = n27644 & n27645;
  assign n27647 = ~n27644 & ~n27645;
  assign n27648 = ~n27646 & ~n27647;
  assign n27649 = n9331 & n26063;
  assign n27650 = n8418 & n22315;
  assign n27651 = n8860 & n22309;
  assign n27652 = ~n27650 & ~n27651;
  assign n27653 = ~n27649 & n27652;
  assign n27654 = ~n8421 & n27653;
  assign n27655 = n26604 & n27653;
  assign n27656 = ~n27654 & ~n27655;
  assign n27657 =  a[8]  & ~n27656;
  assign n27658 = ~ a[8]  & n27656;
  assign n27659 = ~n27657 & ~n27658;
  assign n27660 = n27648 & ~n27659;
  assign n27661 = n27648 & ~n27660;
  assign n27662 = ~n27659 & ~n27660;
  assign n27663 = ~n27661 & ~n27662;
  assign n27664 = ~n27482 & ~n27663;
  assign n27665 = ~n27482 & ~n27664;
  assign n27666 = ~n27663 & ~n27664;
  assign n27667 = ~n27665 & ~n27666;
  assign n27668 = ~n27481 & ~n27667;
  assign n27669 = ~n27481 & ~n27668;
  assign n27670 = ~n27667 & ~n27668;
  assign n27671 = ~n27669 & ~n27670;
  assign n27672 = ~n27400 & ~n27406;
  assign n27673 = n27671 & n27672;
  assign n27674 = ~n27671 & ~n27672;
  assign n27675 = ~n27673 & ~n27674;
  assign n27676 = n75 & n14028;
  assign n27677 = n3020 & ~n13438;
  assign n27678 = n3023 & ~n13627;
  assign n27679 = n3028 & n13941;
  assign n27680 = ~n27678 & ~n27679;
  assign n27681 = ~n27677 & n27680;
  assign n27682 = ~n27676 & n27681;
  assign n27683 = ~n27425 & ~n27427;
  assign n27684 = n3839 & ~n27683;
  assign n27685 = ~n3839 & n27683;
  assign n27686 = ~n27684 & ~n27685;
  assign n27687 = ~n27682 & n27686;
  assign n27688 = ~n27682 & ~n27687;
  assign n27689 = n27686 & ~n27687;
  assign n27690 = ~n27688 & ~n27689;
  assign n27691 = ~n27430 & ~n27434;
  assign n27692 = n27690 & n27691;
  assign n27693 = ~n27690 & ~n27691;
  assign n27694 = ~n27692 & ~n27693;
  assign n27695 = ~n27437 & ~n27440;
  assign n27696 = ~n27694 & n27695;
  assign n27697 = n27694 & ~n27695;
  assign n27698 = ~n27696 & ~n27697;
  assign n27699 = n11727 & n27698;
  assign n27700 = n11055 & n27173;
  assign n27701 = n11715 & n27442;
  assign n27702 = ~n27700 & ~n27701;
  assign n27703 = ~n27699 & n27702;
  assign n27704 = ~n11057 & n27703;
  assign n27705 = ~n27451 & ~n27453;
  assign n27706 = n27442 & n27698;
  assign n27707 = ~n27442 & ~n27698;
  assign n27708 = ~n27705 & ~n27707;
  assign n27709 = ~n27706 & n27708;
  assign n27710 = ~n27705 & ~n27709;
  assign n27711 = ~n27706 & ~n27709;
  assign n27712 = ~n27707 & n27711;
  assign n27713 = ~n27710 & ~n27712;
  assign n27714 = n27703 & n27713;
  assign n27715 = ~n27704 & ~n27714;
  assign n27716 =  a[2]  & ~n27715;
  assign n27717 = ~ a[2]  & n27715;
  assign n27718 = ~n27716 & ~n27717;
  assign n27719 = n27675 & ~n27718;
  assign n27720 = ~n27675 & n27718;
  assign n27721 = ~n27719 & ~n27720;
  assign n27722 = ~n27470 & n27721;
  assign n27723 = n27470 & ~n27721;
  assign n27724 = ~n27722 & ~n27723;
  assign n27725 = n27467 & n27724;
  assign n27726 = ~n27467 & ~n27724;
  assign  result[3]  = ~n27725 & ~n27726;
  assign n27728 = ~n27719 & ~n27722;
  assign n27729 = n71 & n27173;
  assign n27730 = n9867 & n26060;
  assign n27731 = n10434 & n26890;
  assign n27732 = ~n27730 & ~n27731;
  assign n27733 = ~n27729 & n27732;
  assign n27734 = n9870 & n27185;
  assign n27735 = n27733 & ~n27734;
  assign n27736 =  a[5]  & ~n27735;
  assign n27737 = ~n27735 & ~n27736;
  assign n27738 =  a[5]  & ~n27736;
  assign n27739 = ~n27737 & ~n27738;
  assign n27740 = ~n27660 & ~n27664;
  assign n27741 = n7983 & n22315;
  assign n27742 = n7291 & n22320;
  assign n27743 = n7632 & n22312;
  assign n27744 = ~n27742 & ~n27743;
  assign n27745 = ~n27741 & n27744;
  assign n27746 = n7294 & n25294;
  assign n27747 = n27745 & ~n27746;
  assign n27748 =  a[11]  & ~n27747;
  assign n27749 = ~n27747 & ~n27748;
  assign n27750 =  a[11]  & ~n27748;
  assign n27751 = ~n27749 & ~n27750;
  assign n27752 = ~n27633 & ~n27637;
  assign n27753 = n6233 & n22332;
  assign n27754 = n5663 & n22338;
  assign n27755 = n5939 & n22335;
  assign n27756 = ~n27754 & ~n27755;
  assign n27757 = ~n27753 & n27756;
  assign n27758 = n5666 & n22542;
  assign n27759 = n27757 & ~n27758;
  assign n27760 =  a[17]  & ~n27759;
  assign n27761 = ~n27759 & ~n27760;
  assign n27762 =  a[17]  & ~n27760;
  assign n27763 = ~n27761 & ~n27762;
  assign n27764 = ~n27606 & ~n27610;
  assign n27765 = n4694 & n22350;
  assign n27766 = n4533 & n22356;
  assign n27767 = n4604 & n22353;
  assign n27768 = ~n27766 & ~n27767;
  assign n27769 = ~n27765 & n27768;
  assign n27770 = n4536 & n23672;
  assign n27771 = n27769 & ~n27770;
  assign n27772 =  a[23]  & ~n27771;
  assign n27773 = ~n27771 & ~n27772;
  assign n27774 =  a[23]  & ~n27772;
  assign n27775 = ~n27773 & ~n27774;
  assign n27776 = ~n27579 & ~n27583;
  assign n27777 = ~n27562 & ~n27565;
  assign n27778 = ~n27543 & ~n27547;
  assign n27779 = n1423 & n2093;
  assign n27780 = n3544 & n27779;
  assign n27781 = n1575 & n27780;
  assign n27782 = ~n111 & n27781;
  assign n27783 = ~n400 & n27782;
  assign n27784 = ~n226 & n27783;
  assign n27785 = ~n206 & n27784;
  assign n27786 = ~n490 & n27785;
  assign n27787 = ~n165 & n27786;
  assign n27788 = ~n791 & n27787;
  assign n27789 = ~n886 & n27788;
  assign n27790 = n1140 & n2092;
  assign n27791 = n1681 & n27790;
  assign n27792 = n1240 & n27791;
  assign n27793 = n526 & n27792;
  assign n27794 = n3040 & n27793;
  assign n27795 = n1709 & n27794;
  assign n27796 = n3127 & n27795;
  assign n27797 = n4388 & n27796;
  assign n27798 = n2012 & n27797;
  assign n27799 = n27789 & n27798;
  assign n27800 = n120 & n27799;
  assign n27801 = n978 & n27800;
  assign n27802 = n570 & n27801;
  assign n27803 = ~n330 & n27802;
  assign n27804 = ~n602 & n27803;
  assign n27805 = ~n107 & n27804;
  assign n27806 = ~n245 & n27805;
  assign n27807 = ~n429 & n27806;
  assign n27808 = n3020 & n22377;
  assign n27809 = n3028 & n22380;
  assign n27810 = n3023 & n22384;
  assign n27811 = n75 & ~n22834;
  assign n27812 = ~n27810 & ~n27811;
  assign n27813 = ~n27809 & n27812;
  assign n27814 = ~n27808 & n27813;
  assign n27815 = ~n27807 & ~n27814;
  assign n27816 = ~n27807 & ~n27815;
  assign n27817 = ~n27814 & ~n27815;
  assign n27818 = ~n27816 & ~n27817;
  assign n27819 = ~n27778 & ~n27818;
  assign n27820 = ~n27778 & ~n27819;
  assign n27821 = ~n27818 & ~n27819;
  assign n27822 = ~n27820 & ~n27821;
  assign n27823 = n3457 & n22368;
  assign n27824 = n3542 & n22374;
  assign n27825 = n3606 & n22371;
  assign n27826 = ~n27824 & ~n27825;
  assign n27827 = ~n27823 & n27826;
  assign n27828 = ~n3368 & n27827;
  assign n27829 = ~n23006 & n27827;
  assign n27830 = ~n27828 & ~n27829;
  assign n27831 =  a[29]  & ~n27830;
  assign n27832 = ~ a[29]  & n27830;
  assign n27833 = ~n27831 & ~n27832;
  assign n27834 = ~n27822 & ~n27833;
  assign n27835 = n27822 & n27833;
  assign n27836 = ~n27834 & ~n27835;
  assign n27837 = ~n27777 & n27836;
  assign n27838 = n27777 & ~n27836;
  assign n27839 = ~n27837 & ~n27838;
  assign n27840 = n3884 & n22359;
  assign n27841 = n3967 & n22365;
  assign n27842 = n4046 & n22362;
  assign n27843 = ~n27841 & ~n27842;
  assign n27844 = ~n27840 & n27843;
  assign n27845 = ~n4050 & n27844;
  assign n27846 = ~n23368 & n27844;
  assign n27847 = ~n27845 & ~n27846;
  assign n27848 =  a[26]  & ~n27847;
  assign n27849 = ~ a[26]  & n27847;
  assign n27850 = ~n27848 & ~n27849;
  assign n27851 = n27839 & ~n27850;
  assign n27852 = n27839 & ~n27851;
  assign n27853 = ~n27850 & ~n27851;
  assign n27854 = ~n27852 & ~n27853;
  assign n27855 = ~n27776 & ~n27854;
  assign n27856 = ~n27776 & ~n27855;
  assign n27857 = ~n27854 & ~n27855;
  assign n27858 = ~n27856 & ~n27857;
  assign n27859 = ~n27775 & ~n27858;
  assign n27860 = ~n27775 & ~n27859;
  assign n27861 = ~n27858 & ~n27859;
  assign n27862 = ~n27860 & ~n27861;
  assign n27863 = ~n27587 & ~n27593;
  assign n27864 = n27862 & n27863;
  assign n27865 = ~n27862 & ~n27863;
  assign n27866 = ~n27864 & ~n27865;
  assign n27867 = n5496 & n22341;
  assign n27868 = n4935 & n22347;
  assign n27869 = n5407 & n22344;
  assign n27870 = ~n27868 & ~n27869;
  assign n27871 = ~n27867 & n27870;
  assign n27872 = ~n4938 & n27871;
  assign n27873 = ~n24142 & n27871;
  assign n27874 = ~n27872 & ~n27873;
  assign n27875 =  a[20]  & ~n27874;
  assign n27876 = ~ a[20]  & n27874;
  assign n27877 = ~n27875 & ~n27876;
  assign n27878 = n27866 & ~n27877;
  assign n27879 = n27866 & ~n27878;
  assign n27880 = ~n27877 & ~n27878;
  assign n27881 = ~n27879 & ~n27880;
  assign n27882 = ~n27764 & ~n27881;
  assign n27883 = ~n27764 & ~n27882;
  assign n27884 = ~n27881 & ~n27882;
  assign n27885 = ~n27883 & ~n27884;
  assign n27886 = ~n27763 & ~n27885;
  assign n27887 = ~n27763 & ~n27886;
  assign n27888 = ~n27885 & ~n27886;
  assign n27889 = ~n27887 & ~n27888;
  assign n27890 = ~n27614 & ~n27620;
  assign n27891 = n27889 & n27890;
  assign n27892 = ~n27889 & ~n27890;
  assign n27893 = ~n27891 & ~n27892;
  assign n27894 = n7101 & n22323;
  assign n27895 = n6402 & n22329;
  assign n27896 = n6951 & n22326;
  assign n27897 = ~n27895 & ~n27896;
  assign n27898 = ~n27894 & n27897;
  assign n27899 = ~n6397 & n27898;
  assign n27900 = ~n24599 & n27898;
  assign n27901 = ~n27899 & ~n27900;
  assign n27902 =  a[14]  & ~n27901;
  assign n27903 = ~ a[14]  & n27901;
  assign n27904 = ~n27902 & ~n27903;
  assign n27905 = n27893 & ~n27904;
  assign n27906 = n27893 & ~n27905;
  assign n27907 = ~n27904 & ~n27905;
  assign n27908 = ~n27906 & ~n27907;
  assign n27909 = ~n27752 & ~n27908;
  assign n27910 = ~n27752 & ~n27909;
  assign n27911 = ~n27908 & ~n27909;
  assign n27912 = ~n27910 & ~n27911;
  assign n27913 = ~n27751 & ~n27912;
  assign n27914 = ~n27751 & ~n27913;
  assign n27915 = ~n27912 & ~n27913;
  assign n27916 = ~n27914 & ~n27915;
  assign n27917 = ~n27641 & ~n27647;
  assign n27918 = n27916 & n27917;
  assign n27919 = ~n27916 & ~n27917;
  assign n27920 = ~n27918 & ~n27919;
  assign n27921 = n9331 & n26066;
  assign n27922 = n8418 & n22309;
  assign n27923 = n8860 & n26063;
  assign n27924 = ~n27922 & ~n27923;
  assign n27925 = ~n27921 & n27924;
  assign n27926 = ~n8421 & n27925;
  assign n27927 = n26624 & n27925;
  assign n27928 = ~n27926 & ~n27927;
  assign n27929 =  a[8]  & ~n27928;
  assign n27930 = ~ a[8]  & n27928;
  assign n27931 = ~n27929 & ~n27930;
  assign n27932 = n27920 & ~n27931;
  assign n27933 = n27920 & ~n27932;
  assign n27934 = ~n27931 & ~n27932;
  assign n27935 = ~n27933 & ~n27934;
  assign n27936 = ~n27740 & ~n27935;
  assign n27937 = ~n27740 & ~n27936;
  assign n27938 = ~n27935 & ~n27936;
  assign n27939 = ~n27937 & ~n27938;
  assign n27940 = ~n27739 & ~n27939;
  assign n27941 = ~n27739 & ~n27940;
  assign n27942 = ~n27939 & ~n27940;
  assign n27943 = ~n27941 & ~n27942;
  assign n27944 = ~n27668 & ~n27674;
  assign n27945 = n27943 & n27944;
  assign n27946 = ~n27943 & ~n27944;
  assign n27947 = ~n27945 & ~n27946;
  assign n27948 = n75 & ~n13951;
  assign n27949 = ~n3020 & ~n3028;
  assign n27950 = ~n13438 & ~n27949;
  assign n27951 = n3023 & n13941;
  assign n27952 = ~n27950 & ~n27951;
  assign n27953 = ~n27948 & n27952;
  assign n27954 = n3839 & n27953;
  assign n27955 = ~n3839 & ~n27953;
  assign n27956 = ~n27954 & ~n27955;
  assign n27957 = ~n27684 & ~n27687;
  assign n27958 = n27956 & n27957;
  assign n27959 = ~n27956 & ~n27957;
  assign n27960 = ~n27958 & ~n27959;
  assign n27961 = ~n27693 & ~n27697;
  assign n27962 = ~n27960 & n27961;
  assign n27963 = n27960 & ~n27961;
  assign n27964 = ~n27962 & ~n27963;
  assign n27965 = n11727 & n27964;
  assign n27966 = n11055 & n27442;
  assign n27967 = n11715 & n27698;
  assign n27968 = ~n27966 & ~n27967;
  assign n27969 = ~n27965 & n27968;
  assign n27970 = ~n11057 & n27969;
  assign n27971 = ~n27698 & ~n27964;
  assign n27972 = n27698 & n27964;
  assign n27973 = ~n27971 & ~n27972;
  assign n27974 = ~n27711 & n27973;
  assign n27975 = n27711 & ~n27973;
  assign n27976 = ~n27974 & ~n27975;
  assign n27977 = n27969 & ~n27976;
  assign n27978 = ~n27970 & ~n27977;
  assign n27979 =  a[2]  & ~n27978;
  assign n27980 = ~ a[2]  & n27978;
  assign n27981 = ~n27979 & ~n27980;
  assign n27982 = n27947 & ~n27981;
  assign n27983 = ~n27947 & n27981;
  assign n27984 = ~n27982 & ~n27983;
  assign n27985 = ~n27728 & n27984;
  assign n27986 = n27728 & ~n27984;
  assign n27987 = ~n27985 & ~n27986;
  assign n27988 = n27725 & n27987;
  assign n27989 = ~n27725 & ~n27987;
  assign  result[4]  = ~n27988 & ~n27989;
  assign n27991 = ~n27982 & ~n27985;
  assign n27992 = n71 & n27442;
  assign n27993 = n9867 & n26890;
  assign n27994 = n10434 & n27173;
  assign n27995 = ~n27993 & ~n27994;
  assign n27996 = ~n27992 & n27995;
  assign n27997 = n9870 & n27455;
  assign n27998 = n27996 & ~n27997;
  assign n27999 =  a[5]  & ~n27998;
  assign n28000 = ~n27998 & ~n27999;
  assign n28001 =  a[5]  & ~n27999;
  assign n28002 = ~n28000 & ~n28001;
  assign n28003 = ~n27932 & ~n27936;
  assign n28004 = n7983 & n22309;
  assign n28005 = n7291 & n22312;
  assign n28006 = n7632 & n22315;
  assign n28007 = ~n28005 & ~n28006;
  assign n28008 = ~n28004 & n28007;
  assign n28009 = n7294 & ~n22529;
  assign n28010 = n28008 & ~n28009;
  assign n28011 =  a[11]  & ~n28010;
  assign n28012 = ~n28010 & ~n28011;
  assign n28013 =  a[11]  & ~n28011;
  assign n28014 = ~n28012 & ~n28013;
  assign n28015 = ~n27905 & ~n27909;
  assign n28016 = n6233 & n22329;
  assign n28017 = n5663 & n22335;
  assign n28018 = n5939 & n22332;
  assign n28019 = ~n28017 & ~n28018;
  assign n28020 = ~n28016 & n28019;
  assign n28021 = n5666 & ~n24633;
  assign n28022 = n28020 & ~n28021;
  assign n28023 =  a[17]  & ~n28022;
  assign n28024 = ~n28022 & ~n28023;
  assign n28025 =  a[17]  & ~n28023;
  assign n28026 = ~n28024 & ~n28025;
  assign n28027 = ~n27878 & ~n27882;
  assign n28028 = n4694 & n22347;
  assign n28029 = n4533 & n22353;
  assign n28030 = n4604 & n22350;
  assign n28031 = ~n28029 & ~n28030;
  assign n28032 = ~n28028 & n28031;
  assign n28033 = n4536 & ~n23659;
  assign n28034 = n28032 & ~n28033;
  assign n28035 =  a[23]  & ~n28034;
  assign n28036 = ~n28034 & ~n28035;
  assign n28037 =  a[23]  & ~n28035;
  assign n28038 = ~n28036 & ~n28037;
  assign n28039 = ~n27851 & ~n27855;
  assign n28040 = ~n27834 & ~n27837;
  assign n28041 = ~n27815 & ~n27819;
  assign n28042 = n207 & n3587;
  assign n28043 = n690 & n28042;
  assign n28044 = n12409 & n28043;
  assign n28045 = n15970 & n28044;
  assign n28046 = n3644 & n28045;
  assign n28047 = n5286 & n28046;
  assign n28048 = n1046 & n28047;
  assign n28049 = ~n469 & n28048;
  assign n28050 = ~n111 & n28049;
  assign n28051 = ~n242 & n28050;
  assign n28052 = ~n171 & n28051;
  assign n28053 = ~n601 & n28052;
  assign n28054 = ~n375 & n28053;
  assign n28055 = ~n493 & n28054;
  assign n28056 = ~n161 & n28055;
  assign n28057 = ~n251 & n28056;
  assign n28058 = ~n158 & n28057;
  assign n28059 = ~n222 & n28058;
  assign n28060 = n3020 & n22374;
  assign n28061 = n3028 & n22377;
  assign n28062 = n3023 & n22380;
  assign n28063 = n75 & n22569;
  assign n28064 = ~n28062 & ~n28063;
  assign n28065 = ~n28061 & n28064;
  assign n28066 = ~n28060 & n28065;
  assign n28067 = ~n28059 & ~n28066;
  assign n28068 = ~n28059 & ~n28067;
  assign n28069 = ~n28066 & ~n28067;
  assign n28070 = ~n28068 & ~n28069;
  assign n28071 = ~n28041 & ~n28070;
  assign n28072 = ~n28041 & ~n28071;
  assign n28073 = ~n28070 & ~n28071;
  assign n28074 = ~n28072 & ~n28073;
  assign n28075 = n3457 & n22365;
  assign n28076 = n3542 & n22371;
  assign n28077 = n3606 & n22368;
  assign n28078 = ~n28076 & ~n28077;
  assign n28079 = ~n28075 & n28078;
  assign n28080 = ~n3368 & n28079;
  assign n28081 = n22993 & n28079;
  assign n28082 = ~n28080 & ~n28081;
  assign n28083 =  a[29]  & ~n28082;
  assign n28084 = ~ a[29]  & n28082;
  assign n28085 = ~n28083 & ~n28084;
  assign n28086 = ~n28074 & ~n28085;
  assign n28087 = n28074 & n28085;
  assign n28088 = ~n28086 & ~n28087;
  assign n28089 = ~n28040 & n28088;
  assign n28090 = n28040 & ~n28088;
  assign n28091 = ~n28089 & ~n28090;
  assign n28092 = n3884 & n22356;
  assign n28093 = n3967 & n22362;
  assign n28094 = n4046 & n22359;
  assign n28095 = ~n28093 & ~n28094;
  assign n28096 = ~n28092 & n28095;
  assign n28097 = ~n4050 & n28096;
  assign n28098 = n23345 & n28096;
  assign n28099 = ~n28097 & ~n28098;
  assign n28100 =  a[26]  & ~n28099;
  assign n28101 = ~ a[26]  & n28099;
  assign n28102 = ~n28100 & ~n28101;
  assign n28103 = n28091 & ~n28102;
  assign n28104 = n28091 & ~n28103;
  assign n28105 = ~n28102 & ~n28103;
  assign n28106 = ~n28104 & ~n28105;
  assign n28107 = ~n28039 & ~n28106;
  assign n28108 = ~n28039 & ~n28107;
  assign n28109 = ~n28106 & ~n28107;
  assign n28110 = ~n28108 & ~n28109;
  assign n28111 = ~n28038 & ~n28110;
  assign n28112 = ~n28038 & ~n28111;
  assign n28113 = ~n28110 & ~n28111;
  assign n28114 = ~n28112 & ~n28113;
  assign n28115 = ~n27859 & ~n27865;
  assign n28116 = n28114 & n28115;
  assign n28117 = ~n28114 & ~n28115;
  assign n28118 = ~n28116 & ~n28117;
  assign n28119 = n5496 & n22338;
  assign n28120 = n4935 & n22344;
  assign n28121 = n5407 & n22341;
  assign n28122 = ~n28120 & ~n28121;
  assign n28123 = ~n28119 & n28122;
  assign n28124 = ~n4938 & n28123;
  assign n28125 = n24188 & n28123;
  assign n28126 = ~n28124 & ~n28125;
  assign n28127 =  a[20]  & ~n28126;
  assign n28128 = ~ a[20]  & n28126;
  assign n28129 = ~n28127 & ~n28128;
  assign n28130 = n28118 & ~n28129;
  assign n28131 = n28118 & ~n28130;
  assign n28132 = ~n28129 & ~n28130;
  assign n28133 = ~n28131 & ~n28132;
  assign n28134 = ~n28027 & ~n28133;
  assign n28135 = ~n28027 & ~n28134;
  assign n28136 = ~n28133 & ~n28134;
  assign n28137 = ~n28135 & ~n28136;
  assign n28138 = ~n28026 & ~n28137;
  assign n28139 = ~n28026 & ~n28138;
  assign n28140 = ~n28137 & ~n28138;
  assign n28141 = ~n28139 & ~n28140;
  assign n28142 = ~n27886 & ~n27892;
  assign n28143 = n28141 & n28142;
  assign n28144 = ~n28141 & ~n28142;
  assign n28145 = ~n28143 & ~n28144;
  assign n28146 = n7101 & n22320;
  assign n28147 = n6402 & n22326;
  assign n28148 = n6951 & n22323;
  assign n28149 = ~n28147 & ~n28148;
  assign n28150 = ~n28146 & n28149;
  assign n28151 = ~n6397 & n28150;
  assign n28152 = n25270 & n28150;
  assign n28153 = ~n28151 & ~n28152;
  assign n28154 =  a[14]  & ~n28153;
  assign n28155 = ~ a[14]  & n28153;
  assign n28156 = ~n28154 & ~n28155;
  assign n28157 = n28145 & ~n28156;
  assign n28158 = n28145 & ~n28157;
  assign n28159 = ~n28156 & ~n28157;
  assign n28160 = ~n28158 & ~n28159;
  assign n28161 = ~n28015 & ~n28160;
  assign n28162 = ~n28015 & ~n28161;
  assign n28163 = ~n28160 & ~n28161;
  assign n28164 = ~n28162 & ~n28163;
  assign n28165 = ~n28014 & ~n28164;
  assign n28166 = ~n28014 & ~n28165;
  assign n28167 = ~n28164 & ~n28165;
  assign n28168 = ~n28166 & ~n28167;
  assign n28169 = ~n27913 & ~n27919;
  assign n28170 = n28168 & n28169;
  assign n28171 = ~n28168 & ~n28169;
  assign n28172 = ~n28170 & ~n28171;
  assign n28173 = n9331 & n26060;
  assign n28174 = n8418 & n26063;
  assign n28175 = n8860 & n26066;
  assign n28176 = ~n28174 & ~n28175;
  assign n28177 = ~n28173 & n28176;
  assign n28178 = ~n8421 & n28177;
  assign n28179 = n26088 & n28177;
  assign n28180 = ~n28178 & ~n28179;
  assign n28181 =  a[8]  & ~n28180;
  assign n28182 = ~ a[8]  & n28180;
  assign n28183 = ~n28181 & ~n28182;
  assign n28184 = n28172 & ~n28183;
  assign n28185 = n28172 & ~n28184;
  assign n28186 = ~n28183 & ~n28184;
  assign n28187 = ~n28185 & ~n28186;
  assign n28188 = ~n28003 & ~n28187;
  assign n28189 = ~n28003 & ~n28188;
  assign n28190 = ~n28187 & ~n28188;
  assign n28191 = ~n28189 & ~n28190;
  assign n28192 = ~n28002 & ~n28191;
  assign n28193 = ~n28002 & ~n28192;
  assign n28194 = ~n28191 & ~n28192;
  assign n28195 = ~n28193 & ~n28194;
  assign n28196 = ~n27940 & ~n27946;
  assign n28197 = n28195 & n28196;
  assign n28198 = ~n28195 & ~n28196;
  assign n28199 = ~n28197 & ~n28198;
  assign n28200 = ~n27959 & ~n27963;
  assign n28201 = ~ a[31]  & n97;
  assign n28202 = ~n13438 & ~n28201;
  assign n28203 = n27954 & ~n28202;
  assign n28204 = ~n27954 & n28202;
  assign n28205 = ~n28203 & ~n28204;
  assign n28206 = n28200 & ~n28205;
  assign n28207 = ~n28200 & n28205;
  assign n28208 = ~n28206 & ~n28207;
  assign n28209 = n11727 & ~n28208;
  assign n28210 = n11055 & n27698;
  assign n28211 = n11715 & n27964;
  assign n28212 = ~n28210 & ~n28211;
  assign n28213 = ~n28209 & n28212;
  assign n28214 = ~n11057 & n28213;
  assign n28215 = ~n27972 & ~n27974;
  assign n28216 = n27964 & ~n28208;
  assign n28217 = ~n27964 & n28208;
  assign n28218 = ~n28215 & ~n28217;
  assign n28219 = ~n28216 & n28218;
  assign n28220 = ~n28215 & ~n28219;
  assign n28221 = ~n28216 & ~n28219;
  assign n28222 = ~n28217 & n28221;
  assign n28223 = ~n28220 & ~n28222;
  assign n28224 = n28213 & n28223;
  assign n28225 = ~n28214 & ~n28224;
  assign n28226 =  a[2]  & ~n28225;
  assign n28227 = ~ a[2]  & n28225;
  assign n28228 = ~n28226 & ~n28227;
  assign n28229 = n28199 & ~n28228;
  assign n28230 = ~n28199 & n28228;
  assign n28231 = ~n28229 & ~n28230;
  assign n28232 = ~n27991 & n28231;
  assign n28233 = n27991 & ~n28231;
  assign n28234 = ~n28232 & ~n28233;
  assign n28235 = n27988 & n28234;
  assign n28236 = ~n27988 & ~n28234;
  assign  result[5]  = ~n28235 & ~n28236;
  assign n28238 = n71 & n27698;
  assign n28239 = n9867 & n27173;
  assign n28240 = n10434 & n27442;
  assign n28241 = ~n28239 & ~n28240;
  assign n28242 = ~n28238 & n28241;
  assign n28243 = n9870 & ~n27713;
  assign n28244 = n28242 & ~n28243;
  assign n28245 =  a[5]  & ~n28244;
  assign n28246 = ~n28244 & ~n28245;
  assign n28247 =  a[5]  & ~n28245;
  assign n28248 = ~n28246 & ~n28247;
  assign n28249 = ~n28184 & ~n28188;
  assign n28250 = n7983 & n26063;
  assign n28251 = n7291 & n22315;
  assign n28252 = n7632 & n22309;
  assign n28253 = ~n28251 & ~n28252;
  assign n28254 = ~n28250 & n28253;
  assign n28255 = n7294 & ~n26604;
  assign n28256 = n28254 & ~n28255;
  assign n28257 =  a[11]  & ~n28256;
  assign n28258 = ~n28256 & ~n28257;
  assign n28259 =  a[11]  & ~n28257;
  assign n28260 = ~n28258 & ~n28259;
  assign n28261 = ~n28157 & ~n28161;
  assign n28262 = n6233 & n22326;
  assign n28263 = n5663 & n22332;
  assign n28264 = n5939 & n22329;
  assign n28265 = ~n28263 & ~n28264;
  assign n28266 = ~n28262 & n28265;
  assign n28267 = n5666 & ~n24616;
  assign n28268 = n28266 & ~n28267;
  assign n28269 =  a[17]  & ~n28268;
  assign n28270 = ~n28268 & ~n28269;
  assign n28271 =  a[17]  & ~n28269;
  assign n28272 = ~n28270 & ~n28271;
  assign n28273 = ~n28130 & ~n28134;
  assign n28274 = n4694 & n22344;
  assign n28275 = n4533 & n22350;
  assign n28276 = n4604 & n22347;
  assign n28277 = ~n28275 & ~n28276;
  assign n28278 = ~n28274 & n28277;
  assign n28279 = n4536 & ~n23642;
  assign n28280 = n28278 & ~n28279;
  assign n28281 =  a[23]  & ~n28280;
  assign n28282 = ~n28280 & ~n28281;
  assign n28283 =  a[23]  & ~n28281;
  assign n28284 = ~n28282 & ~n28283;
  assign n28285 = ~n28103 & ~n28107;
  assign n28286 = ~n28086 & ~n28089;
  assign n28287 = ~n28067 & ~n28071;
  assign n28288 = n1550 & n1693;
  assign n28289 = ~n169 & n28288;
  assign n28290 = ~n228 & n28289;
  assign n28291 = ~n191 & n28290;
  assign n28292 = ~n567 & n28291;
  assign n28293 = ~n325 & n28292;
  assign n28294 = ~n158 & n28293;
  assign n28295 = n297 & n27522;
  assign n28296 = n437 & n28295;
  assign n28297 = n3040 & n28296;
  assign n28298 = n28294 & n28297;
  assign n28299 = n14565 & n28298;
  assign n28300 = n5013 & n28299;
  assign n28301 = n15047 & n28300;
  assign n28302 = n507 & n28301;
  assign n28303 = n978 & n28302;
  assign n28304 = n227 & n28303;
  assign n28305 = n2405 & n28304;
  assign n28306 = n116 & n28305;
  assign n28307 = ~n656 & n28306;
  assign n28308 = ~n246 & n28307;
  assign n28309 = ~n372 & n28308;
  assign n28310 = ~n657 & n28309;
  assign n28311 = ~n712 & n28310;
  assign n28312 = ~n95 & n28311;
  assign n28313 = ~n886 & n28312;
  assign n28314 = ~n428 & n28313;
  assign n28315 = n3020 & n22371;
  assign n28316 = n3028 & n22374;
  assign n28317 = n3023 & n22377;
  assign n28318 = n75 & n23025;
  assign n28319 = ~n28317 & ~n28318;
  assign n28320 = ~n28316 & n28319;
  assign n28321 = ~n28315 & n28320;
  assign n28322 = ~n28314 & ~n28321;
  assign n28323 = ~n28314 & ~n28322;
  assign n28324 = ~n28321 & ~n28322;
  assign n28325 = ~n28323 & ~n28324;
  assign n28326 = ~n28287 & ~n28325;
  assign n28327 = ~n28287 & ~n28326;
  assign n28328 = ~n28325 & ~n28326;
  assign n28329 = ~n28327 & ~n28328;
  assign n28330 = n3457 & n22362;
  assign n28331 = n3542 & n22368;
  assign n28332 = n3606 & n22365;
  assign n28333 = ~n28331 & ~n28332;
  assign n28334 = ~n28330 & n28333;
  assign n28335 = ~n3368 & n28334;
  assign n28336 = n23320 & n28334;
  assign n28337 = ~n28335 & ~n28336;
  assign n28338 =  a[29]  & ~n28337;
  assign n28339 = ~ a[29]  & n28337;
  assign n28340 = ~n28338 & ~n28339;
  assign n28341 = ~n28329 & ~n28340;
  assign n28342 = n28329 & n28340;
  assign n28343 = ~n28341 & ~n28342;
  assign n28344 = ~n28286 & n28343;
  assign n28345 = n28286 & ~n28343;
  assign n28346 = ~n28344 & ~n28345;
  assign n28347 = n3884 & n22353;
  assign n28348 = n3967 & n22359;
  assign n28349 = n4046 & n22356;
  assign n28350 = ~n28348 & ~n28349;
  assign n28351 = ~n28347 & n28350;
  assign n28352 = ~n4050 & n28351;
  assign n28353 = n22556 & n28351;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 =  a[26]  & ~n28354;
  assign n28356 = ~ a[26]  & n28354;
  assign n28357 = ~n28355 & ~n28356;
  assign n28358 = n28346 & ~n28357;
  assign n28359 = ~n28346 & n28357;
  assign n28360 = ~n28358 & ~n28359;
  assign n28361 = ~n28285 & n28360;
  assign n28362 = n28285 & ~n28360;
  assign n28363 = ~n28361 & ~n28362;
  assign n28364 = ~n28284 & n28363;
  assign n28365 = ~n28284 & ~n28364;
  assign n28366 = n28363 & ~n28364;
  assign n28367 = ~n28365 & ~n28366;
  assign n28368 = ~n28111 & ~n28117;
  assign n28369 = n28367 & n28368;
  assign n28370 = ~n28367 & ~n28368;
  assign n28371 = ~n28369 & ~n28370;
  assign n28372 = n5496 & n22335;
  assign n28373 = n4935 & n22341;
  assign n28374 = n5407 & n22338;
  assign n28375 = ~n28373 & ~n28374;
  assign n28376 = ~n28372 & n28375;
  assign n28377 = ~n4938 & n28376;
  assign n28378 = n24167 & n28376;
  assign n28379 = ~n28377 & ~n28378;
  assign n28380 =  a[20]  & ~n28379;
  assign n28381 = ~ a[20]  & n28379;
  assign n28382 = ~n28380 & ~n28381;
  assign n28383 = n28371 & ~n28382;
  assign n28384 = ~n28371 & n28382;
  assign n28385 = ~n28383 & ~n28384;
  assign n28386 = ~n28273 & n28385;
  assign n28387 = n28273 & ~n28385;
  assign n28388 = ~n28386 & ~n28387;
  assign n28389 = ~n28272 & n28388;
  assign n28390 = ~n28272 & ~n28389;
  assign n28391 = n28388 & ~n28389;
  assign n28392 = ~n28390 & ~n28391;
  assign n28393 = ~n28138 & ~n28144;
  assign n28394 = n28392 & n28393;
  assign n28395 = ~n28392 & ~n28393;
  assign n28396 = ~n28394 & ~n28395;
  assign n28397 = n7101 & n22312;
  assign n28398 = n6402 & n22323;
  assign n28399 = n6951 & n22320;
  assign n28400 = ~n28398 & ~n28399;
  assign n28401 = ~n28397 & n28400;
  assign n28402 = ~n6397 & n28401;
  assign n28403 = n25315 & n28401;
  assign n28404 = ~n28402 & ~n28403;
  assign n28405 =  a[14]  & ~n28404;
  assign n28406 = ~ a[14]  & n28404;
  assign n28407 = ~n28405 & ~n28406;
  assign n28408 = n28396 & ~n28407;
  assign n28409 = ~n28396 & n28407;
  assign n28410 = ~n28408 & ~n28409;
  assign n28411 = ~n28261 & n28410;
  assign n28412 = n28261 & ~n28410;
  assign n28413 = ~n28411 & ~n28412;
  assign n28414 = ~n28260 & n28413;
  assign n28415 = ~n28260 & ~n28414;
  assign n28416 = n28413 & ~n28414;
  assign n28417 = ~n28415 & ~n28416;
  assign n28418 = ~n28165 & ~n28171;
  assign n28419 = n28417 & n28418;
  assign n28420 = ~n28417 & ~n28418;
  assign n28421 = ~n28419 & ~n28420;
  assign n28422 = n9331 & n26890;
  assign n28423 = n8418 & n26066;
  assign n28424 = n8860 & n26060;
  assign n28425 = ~n28423 & ~n28424;
  assign n28426 = ~n28422 & n28425;
  assign n28427 = ~n8421 & n28426;
  assign n28428 = n26904 & n28426;
  assign n28429 = ~n28427 & ~n28428;
  assign n28430 =  a[8]  & ~n28429;
  assign n28431 = ~ a[8]  & n28429;
  assign n28432 = ~n28430 & ~n28431;
  assign n28433 = n28421 & ~n28432;
  assign n28434 = ~n28421 & n28432;
  assign n28435 = ~n28433 & ~n28434;
  assign n28436 = ~n28249 & n28435;
  assign n28437 = n28249 & ~n28435;
  assign n28438 = ~n28436 & ~n28437;
  assign n28439 = ~n28248 & n28438;
  assign n28440 = ~n28248 & ~n28439;
  assign n28441 = n28438 & ~n28439;
  assign n28442 = ~n28440 & ~n28441;
  assign n28443 = ~n20821 & ~n28208;
  assign n28444 = n11055 & n27964;
  assign n28445 = ~n28443 & ~n28444;
  assign n28446 = n11057 & ~n28221;
  assign n28447 = n28445 & ~n28446;
  assign n28448 =  a[2]  & ~n28447;
  assign n28449 =  a[2]  & ~n28448;
  assign n28450 = ~n28447 & ~n28448;
  assign n28451 = ~n28449 & ~n28450;
  assign n28452 = ~n28442 & ~n28451;
  assign n28453 = ~n28442 & ~n28452;
  assign n28454 = ~n28451 & ~n28452;
  assign n28455 = ~n28453 & ~n28454;
  assign n28456 = ~n28192 & ~n28198;
  assign n28457 = n28455 & n28456;
  assign n28458 = ~n28455 & ~n28456;
  assign n28459 = ~n28457 & ~n28458;
  assign n28460 = ~n28229 & ~n28232;
  assign n28461 = ~n28459 & n28460;
  assign n28462 = n28459 & ~n28460;
  assign n28463 = ~n28461 & ~n28462;
  assign n28464 = n28235 & n28463;
  assign n28465 = ~n28235 & ~n28463;
  assign  result[6]  = ~n28464 & ~n28465;
  assign n28467 = ~n28341 & ~n28344;
  assign n28468 = n75 & n23006;
  assign n28469 = n3020 & n22368;
  assign n28470 = n3023 & n22374;
  assign n28471 = n3028 & n22371;
  assign n28472 = ~n28470 & ~n28471;
  assign n28473 = ~n28469 & n28472;
  assign n28474 = ~n28468 & n28473;
  assign n28475 = n2115 & n2423;
  assign n28476 = n6734 & n28475;
  assign n28477 = n13698 & n28476;
  assign n28478 = n2022 & n28477;
  assign n28479 = n12944 & n28478;
  assign n28480 = n1577 & n28479;
  assign n28481 = n3757 & n28480;
  assign n28482 = n1884 & n28481;
  assign n28483 = n1574 & n28482;
  assign n28484 = n3984 & n28483;
  assign n28485 = n2483 & n28484;
  assign n28486 = n1389 & n28485;
  assign n28487 = ~n847 & n28486;
  assign n28488 = ~n619 & n28487;
  assign n28489 = ~n601 & n28488;
  assign n28490 = ~n537 & n28489;
  assign n28491 = ~n157 & n28490;
  assign n28492 = ~n531 & n28491;
  assign n28493 = ~n15031 & ~n28208;
  assign n28494 =  a[2]  & ~n28493;
  assign n28495 = ~ a[2]  & n28493;
  assign n28496 = ~n28494 & ~n28495;
  assign n28497 = ~n28492 & ~n28496;
  assign n28498 = n28492 & n28496;
  assign n28499 = ~n28474 & ~n28498;
  assign n28500 = ~n28497 & n28499;
  assign n28501 = ~n28474 & ~n28500;
  assign n28502 = ~n28497 & ~n28500;
  assign n28503 = ~n28498 & n28502;
  assign n28504 = ~n28501 & ~n28503;
  assign n28505 = ~n28322 & ~n28326;
  assign n28506 = n28504 & n28505;
  assign n28507 = ~n28504 & ~n28505;
  assign n28508 = ~n28506 & ~n28507;
  assign n28509 = n3457 & n22359;
  assign n28510 = n3542 & n22365;
  assign n28511 = n3606 & n22362;
  assign n28512 = ~n28510 & ~n28511;
  assign n28513 = ~n28509 & n28512;
  assign n28514 = ~n3368 & n28513;
  assign n28515 = ~n23368 & n28513;
  assign n28516 = ~n28514 & ~n28515;
  assign n28517 =  a[29]  & ~n28516;
  assign n28518 = ~ a[29]  & n28516;
  assign n28519 = ~n28517 & ~n28518;
  assign n28520 = n28508 & ~n28519;
  assign n28521 = ~n28508 & n28519;
  assign n28522 = ~n28520 & ~n28521;
  assign n28523 = ~n28467 & n28522;
  assign n28524 = n28467 & ~n28522;
  assign n28525 = ~n28523 & ~n28524;
  assign n28526 = n3884 & n22350;
  assign n28527 = n3967 & n22356;
  assign n28528 = n4046 & n22353;
  assign n28529 = ~n28527 & ~n28528;
  assign n28530 = ~n28526 & n28529;
  assign n28531 = n4050 & n23672;
  assign n28532 = n28530 & ~n28531;
  assign n28533 =  a[26]  & ~n28532;
  assign n28534 =  a[26]  & ~n28533;
  assign n28535 = ~n28532 & ~n28533;
  assign n28536 = ~n28534 & ~n28535;
  assign n28537 = n28525 & ~n28536;
  assign n28538 = n28525 & ~n28537;
  assign n28539 = ~n28536 & ~n28537;
  assign n28540 = ~n28538 & ~n28539;
  assign n28541 = ~n28358 & ~n28361;
  assign n28542 = n28540 & n28541;
  assign n28543 = ~n28540 & ~n28541;
  assign n28544 = ~n28542 & ~n28543;
  assign n28545 = n4694 & n22341;
  assign n28546 = n4533 & n22347;
  assign n28547 = n4604 & n22344;
  assign n28548 = ~n28546 & ~n28547;
  assign n28549 = ~n28545 & n28548;
  assign n28550 = n4536 & n24142;
  assign n28551 = n28549 & ~n28550;
  assign n28552 =  a[23]  & ~n28551;
  assign n28553 =  a[23]  & ~n28552;
  assign n28554 = ~n28551 & ~n28552;
  assign n28555 = ~n28553 & ~n28554;
  assign n28556 = n28544 & ~n28555;
  assign n28557 = n28544 & ~n28556;
  assign n28558 = ~n28555 & ~n28556;
  assign n28559 = ~n28557 & ~n28558;
  assign n28560 = ~n28364 & ~n28370;
  assign n28561 = n28559 & n28560;
  assign n28562 = ~n28559 & ~n28560;
  assign n28563 = ~n28561 & ~n28562;
  assign n28564 = n5496 & n22332;
  assign n28565 = n4935 & n22338;
  assign n28566 = n5407 & n22335;
  assign n28567 = ~n28565 & ~n28566;
  assign n28568 = ~n28564 & n28567;
  assign n28569 = n4938 & n22542;
  assign n28570 = n28568 & ~n28569;
  assign n28571 =  a[20]  & ~n28570;
  assign n28572 =  a[20]  & ~n28571;
  assign n28573 = ~n28570 & ~n28571;
  assign n28574 = ~n28572 & ~n28573;
  assign n28575 = n28563 & ~n28574;
  assign n28576 = n28563 & ~n28575;
  assign n28577 = ~n28574 & ~n28575;
  assign n28578 = ~n28576 & ~n28577;
  assign n28579 = ~n28383 & ~n28386;
  assign n28580 = n28578 & n28579;
  assign n28581 = ~n28578 & ~n28579;
  assign n28582 = ~n28580 & ~n28581;
  assign n28583 = n6233 & n22323;
  assign n28584 = n5663 & n22329;
  assign n28585 = n5939 & n22326;
  assign n28586 = ~n28584 & ~n28585;
  assign n28587 = ~n28583 & n28586;
  assign n28588 = n5666 & n24599;
  assign n28589 = n28587 & ~n28588;
  assign n28590 =  a[17]  & ~n28589;
  assign n28591 =  a[17]  & ~n28590;
  assign n28592 = ~n28589 & ~n28590;
  assign n28593 = ~n28591 & ~n28592;
  assign n28594 = n28582 & ~n28593;
  assign n28595 = n28582 & ~n28594;
  assign n28596 = ~n28593 & ~n28594;
  assign n28597 = ~n28595 & ~n28596;
  assign n28598 = ~n28389 & ~n28395;
  assign n28599 = n28597 & n28598;
  assign n28600 = ~n28597 & ~n28598;
  assign n28601 = ~n28599 & ~n28600;
  assign n28602 = n7101 & n22315;
  assign n28603 = n6402 & n22320;
  assign n28604 = n6951 & n22312;
  assign n28605 = ~n28603 & ~n28604;
  assign n28606 = ~n28602 & n28605;
  assign n28607 = n6397 & n25294;
  assign n28608 = n28606 & ~n28607;
  assign n28609 =  a[14]  & ~n28608;
  assign n28610 =  a[14]  & ~n28609;
  assign n28611 = ~n28608 & ~n28609;
  assign n28612 = ~n28610 & ~n28611;
  assign n28613 = n28601 & ~n28612;
  assign n28614 = n28601 & ~n28613;
  assign n28615 = ~n28612 & ~n28613;
  assign n28616 = ~n28614 & ~n28615;
  assign n28617 = ~n28408 & ~n28411;
  assign n28618 = n28616 & n28617;
  assign n28619 = ~n28616 & ~n28617;
  assign n28620 = ~n28618 & ~n28619;
  assign n28621 = n7983 & n26066;
  assign n28622 = n7291 & n22309;
  assign n28623 = n7632 & n26063;
  assign n28624 = ~n28622 & ~n28623;
  assign n28625 = ~n28621 & n28624;
  assign n28626 = n7294 & ~n26624;
  assign n28627 = n28625 & ~n28626;
  assign n28628 =  a[11]  & ~n28627;
  assign n28629 =  a[11]  & ~n28628;
  assign n28630 = ~n28627 & ~n28628;
  assign n28631 = ~n28629 & ~n28630;
  assign n28632 = n28620 & ~n28631;
  assign n28633 = n28620 & ~n28632;
  assign n28634 = ~n28631 & ~n28632;
  assign n28635 = ~n28633 & ~n28634;
  assign n28636 = ~n28414 & ~n28420;
  assign n28637 = n28635 & n28636;
  assign n28638 = ~n28635 & ~n28636;
  assign n28639 = ~n28637 & ~n28638;
  assign n28640 = n9331 & n27173;
  assign n28641 = n8418 & n26060;
  assign n28642 = n8860 & n26890;
  assign n28643 = ~n28641 & ~n28642;
  assign n28644 = ~n28640 & n28643;
  assign n28645 = n8421 & n27185;
  assign n28646 = n28644 & ~n28645;
  assign n28647 =  a[8]  & ~n28646;
  assign n28648 =  a[8]  & ~n28647;
  assign n28649 = ~n28646 & ~n28647;
  assign n28650 = ~n28648 & ~n28649;
  assign n28651 = n28639 & ~n28650;
  assign n28652 = n28639 & ~n28651;
  assign n28653 = ~n28650 & ~n28651;
  assign n28654 = ~n28652 & ~n28653;
  assign n28655 = ~n28433 & ~n28436;
  assign n28656 = n28654 & n28655;
  assign n28657 = ~n28654 & ~n28655;
  assign n28658 = ~n28656 & ~n28657;
  assign n28659 = n71 & n27964;
  assign n28660 = n9867 & n27442;
  assign n28661 = n10434 & n27698;
  assign n28662 = ~n28660 & ~n28661;
  assign n28663 = ~n28659 & n28662;
  assign n28664 = n9870 & n27976;
  assign n28665 = n28663 & ~n28664;
  assign n28666 =  a[5]  & ~n28665;
  assign n28667 =  a[5]  & ~n28666;
  assign n28668 = ~n28665 & ~n28666;
  assign n28669 = ~n28667 & ~n28668;
  assign n28670 = n28658 & ~n28669;
  assign n28671 = n28658 & ~n28670;
  assign n28672 = ~n28669 & ~n28670;
  assign n28673 = ~n28671 & ~n28672;
  assign n28674 = ~n28439 & ~n28452;
  assign n28675 = n28673 & n28674;
  assign n28676 = ~n28673 & ~n28674;
  assign n28677 = ~n28675 & ~n28676;
  assign n28678 = ~n28458 & ~n28462;
  assign n28679 = ~n28677 & n28678;
  assign n28680 = n28677 & ~n28678;
  assign n28681 = ~n28679 & ~n28680;
  assign n28682 = n28464 & n28681;
  assign n28683 = ~n28464 & ~n28681;
  assign  result[7]  = ~n28682 & ~n28683;
  assign n28685 = n720 & n16020;
  assign n28686 = ~n301 & n28685;
  assign n28687 = ~n571 & n28686;
  assign n28688 = ~n886 & n28687;
  assign n28689 = n1347 & n23251;
  assign n28690 = n1424 & n28689;
  assign n28691 = n2410 & n28690;
  assign n28692 = n28688 & n28691;
  assign n28693 = n16067 & n28692;
  assign n28694 = n1313 & n28693;
  assign n28695 = n1782 & n28694;
  assign n28696 = n869 & n28695;
  assign n28697 = n979 & n28696;
  assign n28698 = n399 & n28697;
  assign n28699 = n2583 & n28698;
  assign n28700 = n2088 & n28699;
  assign n28701 = n3163 & n28700;
  assign n28702 = n279 & n28701;
  assign n28703 = ~n121 & n28702;
  assign n28704 = ~n283 & n28703;
  assign n28705 = ~n666 & n28704;
  assign n28706 = ~n363 & n28705;
  assign n28707 = ~n28496 & ~n28706;
  assign n28708 = n28496 & n28706;
  assign n28709 = ~n28502 & ~n28708;
  assign n28710 = ~n28707 & n28709;
  assign n28711 = ~n28502 & ~n28710;
  assign n28712 = ~n28707 & ~n28710;
  assign n28713 = ~n28708 & n28712;
  assign n28714 = ~n28711 & ~n28713;
  assign n28715 = n75 & ~n22993;
  assign n28716 = n3020 & n22365;
  assign n28717 = n3023 & n22371;
  assign n28718 = n3028 & n22368;
  assign n28719 = ~n28717 & ~n28718;
  assign n28720 = ~n28716 & n28719;
  assign n28721 = ~n28715 & n28720;
  assign n28722 = ~n28714 & ~n28721;
  assign n28723 = ~n28714 & ~n28722;
  assign n28724 = ~n28721 & ~n28722;
  assign n28725 = ~n28723 & ~n28724;
  assign n28726 = ~n28507 & ~n28520;
  assign n28727 = n28725 & n28726;
  assign n28728 = ~n28725 & ~n28726;
  assign n28729 = ~n28727 & ~n28728;
  assign n28730 = n3457 & n22356;
  assign n28731 = n3542 & n22362;
  assign n28732 = n3606 & n22359;
  assign n28733 = ~n28731 & ~n28732;
  assign n28734 = ~n28730 & n28733;
  assign n28735 = n3368 & ~n23345;
  assign n28736 = n28734 & ~n28735;
  assign n28737 =  a[29]  & ~n28736;
  assign n28738 =  a[29]  & ~n28737;
  assign n28739 = ~n28736 & ~n28737;
  assign n28740 = ~n28738 & ~n28739;
  assign n28741 = n28729 & ~n28740;
  assign n28742 = n28729 & ~n28741;
  assign n28743 = ~n28740 & ~n28741;
  assign n28744 = ~n28742 & ~n28743;
  assign n28745 = n3884 & n22347;
  assign n28746 = n3967 & n22353;
  assign n28747 = n4046 & n22350;
  assign n28748 = ~n28746 & ~n28747;
  assign n28749 = ~n28745 & n28748;
  assign n28750 = n4050 & ~n23659;
  assign n28751 = n28749 & ~n28750;
  assign n28752 =  a[26]  & ~n28751;
  assign n28753 =  a[26]  & ~n28752;
  assign n28754 = ~n28751 & ~n28752;
  assign n28755 = ~n28753 & ~n28754;
  assign n28756 = ~n28744 & ~n28755;
  assign n28757 = ~n28744 & ~n28756;
  assign n28758 = ~n28755 & ~n28756;
  assign n28759 = ~n28757 & ~n28758;
  assign n28760 = ~n28523 & ~n28537;
  assign n28761 = n28759 & n28760;
  assign n28762 = ~n28759 & ~n28760;
  assign n28763 = ~n28761 & ~n28762;
  assign n28764 = n4694 & n22338;
  assign n28765 = n4533 & n22344;
  assign n28766 = n4604 & n22341;
  assign n28767 = ~n28765 & ~n28766;
  assign n28768 = ~n28764 & n28767;
  assign n28769 = n4536 & ~n24188;
  assign n28770 = n28768 & ~n28769;
  assign n28771 =  a[23]  & ~n28770;
  assign n28772 =  a[23]  & ~n28771;
  assign n28773 = ~n28770 & ~n28771;
  assign n28774 = ~n28772 & ~n28773;
  assign n28775 = n28763 & ~n28774;
  assign n28776 = n28763 & ~n28775;
  assign n28777 = ~n28774 & ~n28775;
  assign n28778 = ~n28776 & ~n28777;
  assign n28779 = ~n28543 & ~n28556;
  assign n28780 = n28778 & n28779;
  assign n28781 = ~n28778 & ~n28779;
  assign n28782 = ~n28780 & ~n28781;
  assign n28783 = n5496 & n22329;
  assign n28784 = n4935 & n22335;
  assign n28785 = n5407 & n22332;
  assign n28786 = ~n28784 & ~n28785;
  assign n28787 = ~n28783 & n28786;
  assign n28788 = n4938 & ~n24633;
  assign n28789 = n28787 & ~n28788;
  assign n28790 =  a[20]  & ~n28789;
  assign n28791 =  a[20]  & ~n28790;
  assign n28792 = ~n28789 & ~n28790;
  assign n28793 = ~n28791 & ~n28792;
  assign n28794 = n28782 & ~n28793;
  assign n28795 = n28782 & ~n28794;
  assign n28796 = ~n28793 & ~n28794;
  assign n28797 = ~n28795 & ~n28796;
  assign n28798 = ~n28562 & ~n28575;
  assign n28799 = n28797 & n28798;
  assign n28800 = ~n28797 & ~n28798;
  assign n28801 = ~n28799 & ~n28800;
  assign n28802 = n6233 & n22320;
  assign n28803 = n5663 & n22326;
  assign n28804 = n5939 & n22323;
  assign n28805 = ~n28803 & ~n28804;
  assign n28806 = ~n28802 & n28805;
  assign n28807 = n5666 & ~n25270;
  assign n28808 = n28806 & ~n28807;
  assign n28809 =  a[17]  & ~n28808;
  assign n28810 =  a[17]  & ~n28809;
  assign n28811 = ~n28808 & ~n28809;
  assign n28812 = ~n28810 & ~n28811;
  assign n28813 = n28801 & ~n28812;
  assign n28814 = n28801 & ~n28813;
  assign n28815 = ~n28812 & ~n28813;
  assign n28816 = ~n28814 & ~n28815;
  assign n28817 = ~n28581 & ~n28594;
  assign n28818 = n28816 & n28817;
  assign n28819 = ~n28816 & ~n28817;
  assign n28820 = ~n28818 & ~n28819;
  assign n28821 = n7101 & n22309;
  assign n28822 = n6402 & n22312;
  assign n28823 = n6951 & n22315;
  assign n28824 = ~n28822 & ~n28823;
  assign n28825 = ~n28821 & n28824;
  assign n28826 = n6397 & ~n22529;
  assign n28827 = n28825 & ~n28826;
  assign n28828 =  a[14]  & ~n28827;
  assign n28829 =  a[14]  & ~n28828;
  assign n28830 = ~n28827 & ~n28828;
  assign n28831 = ~n28829 & ~n28830;
  assign n28832 = n28820 & ~n28831;
  assign n28833 = n28820 & ~n28832;
  assign n28834 = ~n28831 & ~n28832;
  assign n28835 = ~n28833 & ~n28834;
  assign n28836 = ~n28600 & ~n28613;
  assign n28837 = n28835 & n28836;
  assign n28838 = ~n28835 & ~n28836;
  assign n28839 = ~n28837 & ~n28838;
  assign n28840 = n7983 & n26060;
  assign n28841 = n7291 & n26063;
  assign n28842 = n7632 & n26066;
  assign n28843 = ~n28841 & ~n28842;
  assign n28844 = ~n28840 & n28843;
  assign n28845 = n7294 & ~n26088;
  assign n28846 = n28844 & ~n28845;
  assign n28847 =  a[11]  & ~n28846;
  assign n28848 =  a[11]  & ~n28847;
  assign n28849 = ~n28846 & ~n28847;
  assign n28850 = ~n28848 & ~n28849;
  assign n28851 = n28839 & ~n28850;
  assign n28852 = n28839 & ~n28851;
  assign n28853 = ~n28850 & ~n28851;
  assign n28854 = ~n28852 & ~n28853;
  assign n28855 = ~n28619 & ~n28632;
  assign n28856 = n28854 & n28855;
  assign n28857 = ~n28854 & ~n28855;
  assign n28858 = ~n28856 & ~n28857;
  assign n28859 = n9331 & n27442;
  assign n28860 = n8418 & n26890;
  assign n28861 = n8860 & n27173;
  assign n28862 = ~n28860 & ~n28861;
  assign n28863 = ~n28859 & n28862;
  assign n28864 = n8421 & n27455;
  assign n28865 = n28863 & ~n28864;
  assign n28866 =  a[8]  & ~n28865;
  assign n28867 =  a[8]  & ~n28866;
  assign n28868 = ~n28865 & ~n28866;
  assign n28869 = ~n28867 & ~n28868;
  assign n28870 = n28858 & ~n28869;
  assign n28871 = n28858 & ~n28870;
  assign n28872 = ~n28869 & ~n28870;
  assign n28873 = ~n28871 & ~n28872;
  assign n28874 = ~n28638 & ~n28651;
  assign n28875 = n28873 & n28874;
  assign n28876 = ~n28873 & ~n28874;
  assign n28877 = ~n28875 & ~n28876;
  assign n28878 = n71 & ~n28208;
  assign n28879 = n9867 & n27698;
  assign n28880 = n10434 & n27964;
  assign n28881 = ~n28879 & ~n28880;
  assign n28882 = ~n28878 & n28881;
  assign n28883 = n9870 & ~n28223;
  assign n28884 = n28882 & ~n28883;
  assign n28885 =  a[5]  & ~n28884;
  assign n28886 =  a[5]  & ~n28885;
  assign n28887 = ~n28884 & ~n28885;
  assign n28888 = ~n28886 & ~n28887;
  assign n28889 = n28877 & ~n28888;
  assign n28890 = n28877 & ~n28889;
  assign n28891 = ~n28888 & ~n28889;
  assign n28892 = ~n28890 & ~n28891;
  assign n28893 = ~n28657 & ~n28670;
  assign n28894 = n28892 & n28893;
  assign n28895 = ~n28892 & ~n28893;
  assign n28896 = ~n28894 & ~n28895;
  assign n28897 = ~n28676 & ~n28680;
  assign n28898 = ~n28896 & n28897;
  assign n28899 = n28896 & ~n28897;
  assign n28900 = ~n28898 & ~n28899;
  assign n28901 = n28682 & n28900;
  assign n28902 = ~n28682 & ~n28900;
  assign  result[8]  = ~n28901 & ~n28902;
  assign n28904 = n2424 & n15286;
  assign n28905 = n2704 & n28904;
  assign n28906 = n1103 & n28905;
  assign n28907 = n3685 & n28906;
  assign n28908 = n5199 & n28907;
  assign n28909 = n770 & n28908;
  assign n28910 = n415 & n28909;
  assign n28911 = n1182 & n28910;
  assign n28912 = n2443 & n28911;
  assign n28913 = n937 & n28912;
  assign n28914 = n2167 & n28913;
  assign n28915 = ~n276 & n28914;
  assign n28916 = ~n1011 & n28915;
  assign n28917 = ~n255 & n28916;
  assign n28918 = ~n150 & n28917;
  assign n28919 = ~n295 & n28918;
  assign n28920 = ~n28496 & ~n28919;
  assign n28921 = n28496 & n28919;
  assign n28922 = ~n28712 & ~n28921;
  assign n28923 = ~n28920 & n28922;
  assign n28924 = ~n28712 & ~n28923;
  assign n28925 = ~n28920 & ~n28923;
  assign n28926 = ~n28921 & n28925;
  assign n28927 = ~n28924 & ~n28926;
  assign n28928 = n75 & ~n23320;
  assign n28929 = n3020 & n22362;
  assign n28930 = n3023 & n22368;
  assign n28931 = n3028 & n22365;
  assign n28932 = ~n28930 & ~n28931;
  assign n28933 = ~n28929 & n28932;
  assign n28934 = ~n28928 & n28933;
  assign n28935 = ~n28927 & ~n28934;
  assign n28936 = ~n28927 & ~n28935;
  assign n28937 = ~n28934 & ~n28935;
  assign n28938 = ~n28936 & ~n28937;
  assign n28939 = ~n28722 & ~n28728;
  assign n28940 = n28938 & n28939;
  assign n28941 = ~n28938 & ~n28939;
  assign n28942 = ~n28940 & ~n28941;
  assign n28943 = n3457 & n22353;
  assign n28944 = n3542 & n22359;
  assign n28945 = n3606 & n22356;
  assign n28946 = ~n28944 & ~n28945;
  assign n28947 = ~n28943 & n28946;
  assign n28948 = n3368 & ~n22556;
  assign n28949 = n28947 & ~n28948;
  assign n28950 =  a[29]  & ~n28949;
  assign n28951 =  a[29]  & ~n28950;
  assign n28952 = ~n28949 & ~n28950;
  assign n28953 = ~n28951 & ~n28952;
  assign n28954 = n28942 & ~n28953;
  assign n28955 = n28942 & ~n28954;
  assign n28956 = ~n28953 & ~n28954;
  assign n28957 = ~n28955 & ~n28956;
  assign n28958 = n3884 & n22344;
  assign n28959 = n3967 & n22350;
  assign n28960 = n4046 & n22347;
  assign n28961 = ~n28959 & ~n28960;
  assign n28962 = ~n28958 & n28961;
  assign n28963 = n4050 & ~n23642;
  assign n28964 = n28962 & ~n28963;
  assign n28965 =  a[26]  & ~n28964;
  assign n28966 =  a[26]  & ~n28965;
  assign n28967 = ~n28964 & ~n28965;
  assign n28968 = ~n28966 & ~n28967;
  assign n28969 = ~n28957 & ~n28968;
  assign n28970 = ~n28957 & ~n28969;
  assign n28971 = ~n28968 & ~n28969;
  assign n28972 = ~n28970 & ~n28971;
  assign n28973 = ~n28741 & ~n28756;
  assign n28974 = n28972 & n28973;
  assign n28975 = ~n28972 & ~n28973;
  assign n28976 = ~n28974 & ~n28975;
  assign n28977 = n4694 & n22335;
  assign n28978 = n4533 & n22341;
  assign n28979 = n4604 & n22338;
  assign n28980 = ~n28978 & ~n28979;
  assign n28981 = ~n28977 & n28980;
  assign n28982 = n4536 & ~n24167;
  assign n28983 = n28981 & ~n28982;
  assign n28984 =  a[23]  & ~n28983;
  assign n28985 =  a[23]  & ~n28984;
  assign n28986 = ~n28983 & ~n28984;
  assign n28987 = ~n28985 & ~n28986;
  assign n28988 = n28976 & ~n28987;
  assign n28989 = n28976 & ~n28988;
  assign n28990 = ~n28987 & ~n28988;
  assign n28991 = ~n28989 & ~n28990;
  assign n28992 = ~n28762 & ~n28775;
  assign n28993 = n28991 & n28992;
  assign n28994 = ~n28991 & ~n28992;
  assign n28995 = ~n28993 & ~n28994;
  assign n28996 = n5496 & n22326;
  assign n28997 = n4935 & n22332;
  assign n28998 = n5407 & n22329;
  assign n28999 = ~n28997 & ~n28998;
  assign n29000 = ~n28996 & n28999;
  assign n29001 = n4938 & ~n24616;
  assign n29002 = n29000 & ~n29001;
  assign n29003 =  a[20]  & ~n29002;
  assign n29004 =  a[20]  & ~n29003;
  assign n29005 = ~n29002 & ~n29003;
  assign n29006 = ~n29004 & ~n29005;
  assign n29007 = n28995 & ~n29006;
  assign n29008 = n28995 & ~n29007;
  assign n29009 = ~n29006 & ~n29007;
  assign n29010 = ~n29008 & ~n29009;
  assign n29011 = ~n28781 & ~n28794;
  assign n29012 = n29010 & n29011;
  assign n29013 = ~n29010 & ~n29011;
  assign n29014 = ~n29012 & ~n29013;
  assign n29015 = n6233 & n22312;
  assign n29016 = n5663 & n22323;
  assign n29017 = n5939 & n22320;
  assign n29018 = ~n29016 & ~n29017;
  assign n29019 = ~n29015 & n29018;
  assign n29020 = n5666 & ~n25315;
  assign n29021 = n29019 & ~n29020;
  assign n29022 =  a[17]  & ~n29021;
  assign n29023 =  a[17]  & ~n29022;
  assign n29024 = ~n29021 & ~n29022;
  assign n29025 = ~n29023 & ~n29024;
  assign n29026 = n29014 & ~n29025;
  assign n29027 = n29014 & ~n29026;
  assign n29028 = ~n29025 & ~n29026;
  assign n29029 = ~n29027 & ~n29028;
  assign n29030 = ~n28800 & ~n28813;
  assign n29031 = n29029 & n29030;
  assign n29032 = ~n29029 & ~n29030;
  assign n29033 = ~n29031 & ~n29032;
  assign n29034 = n7101 & n26063;
  assign n29035 = n6402 & n22315;
  assign n29036 = n6951 & n22309;
  assign n29037 = ~n29035 & ~n29036;
  assign n29038 = ~n29034 & n29037;
  assign n29039 = n6397 & ~n26604;
  assign n29040 = n29038 & ~n29039;
  assign n29041 =  a[14]  & ~n29040;
  assign n29042 =  a[14]  & ~n29041;
  assign n29043 = ~n29040 & ~n29041;
  assign n29044 = ~n29042 & ~n29043;
  assign n29045 = n29033 & ~n29044;
  assign n29046 = n29033 & ~n29045;
  assign n29047 = ~n29044 & ~n29045;
  assign n29048 = ~n29046 & ~n29047;
  assign n29049 = ~n28819 & ~n28832;
  assign n29050 = n29048 & n29049;
  assign n29051 = ~n29048 & ~n29049;
  assign n29052 = ~n29050 & ~n29051;
  assign n29053 = n7983 & n26890;
  assign n29054 = n7291 & n26066;
  assign n29055 = n7632 & n26060;
  assign n29056 = ~n29054 & ~n29055;
  assign n29057 = ~n29053 & n29056;
  assign n29058 = n7294 & ~n26904;
  assign n29059 = n29057 & ~n29058;
  assign n29060 =  a[11]  & ~n29059;
  assign n29061 =  a[11]  & ~n29060;
  assign n29062 = ~n29059 & ~n29060;
  assign n29063 = ~n29061 & ~n29062;
  assign n29064 = n29052 & ~n29063;
  assign n29065 = n29052 & ~n29064;
  assign n29066 = ~n29063 & ~n29064;
  assign n29067 = ~n29065 & ~n29066;
  assign n29068 = ~n28838 & ~n28851;
  assign n29069 = n29067 & n29068;
  assign n29070 = ~n29067 & ~n29068;
  assign n29071 = ~n29069 & ~n29070;
  assign n29072 = n9331 & n27698;
  assign n29073 = n8418 & n27173;
  assign n29074 = n8860 & n27442;
  assign n29075 = ~n29073 & ~n29074;
  assign n29076 = ~n29072 & n29075;
  assign n29077 = n8421 & ~n27713;
  assign n29078 = n29076 & ~n29077;
  assign n29079 =  a[8]  & ~n29078;
  assign n29080 =  a[8]  & ~n29079;
  assign n29081 = ~n29078 & ~n29079;
  assign n29082 = ~n29080 & ~n29081;
  assign n29083 = n29071 & ~n29082;
  assign n29084 = n29071 & ~n29083;
  assign n29085 = ~n29082 & ~n29083;
  assign n29086 = ~n29084 & ~n29085;
  assign n29087 = ~n28857 & ~n28870;
  assign n29088 = ~n15076 & ~n28208;
  assign n29089 = n9867 & n27964;
  assign n29090 = ~n29088 & ~n29089;
  assign n29091 = ~n9870 & n29090;
  assign n29092 = n28221 & n29090;
  assign n29093 = ~n29091 & ~n29092;
  assign n29094 =  a[5]  & ~n29093;
  assign n29095 = ~ a[5]  & n29093;
  assign n29096 = ~n29094 & ~n29095;
  assign n29097 = ~n29087 & ~n29096;
  assign n29098 = n29087 & n29096;
  assign n29099 = ~n29097 & ~n29098;
  assign n29100 = ~n29086 & n29099;
  assign n29101 = ~n29086 & ~n29100;
  assign n29102 = n29099 & ~n29100;
  assign n29103 = ~n29101 & ~n29102;
  assign n29104 = ~n28876 & ~n28889;
  assign n29105 = n29103 & n29104;
  assign n29106 = ~n29103 & ~n29104;
  assign n29107 = ~n29105 & ~n29106;
  assign n29108 = ~n28895 & ~n28899;
  assign n29109 = ~n29107 & n29108;
  assign n29110 = n29107 & ~n29108;
  assign n29111 = ~n29109 & ~n29110;
  assign n29112 = n28901 & n29111;
  assign n29113 = ~n28901 & ~n29111;
  assign  result[9]  = ~n29112 & ~n29113;
  assign n29115 = ~n29106 & ~n29110;
  assign n29116 = ~n29097 & ~n29100;
  assign n29117 = ~n28935 & ~n28941;
  assign n29118 = n1859 & n4335;
  assign n29119 = n1073 & n29118;
  assign n29120 = n4357 & n29119;
  assign n29121 = n960 & n29120;
  assign n29122 = n526 & n29121;
  assign n29123 = n13826 & n29122;
  assign n29124 = n3057 & n29123;
  assign n29125 = n2467 & n29124;
  assign n29126 = n3886 & n29125;
  assign n29127 = n1761 & n29126;
  assign n29128 = n22748 & n29127;
  assign n29129 = ~n746 & n29128;
  assign n29130 = ~n280 & n29129;
  assign n29131 = ~n119 & n29130;
  assign n29132 = ~n358 & n29131;
  assign n29133 = n28496 & n29132;
  assign n29134 = ~n28496 & ~n29132;
  assign n29135 = ~n29133 & ~n29134;
  assign n29136 = ~n15078 & ~n28208;
  assign n29137 = ~ a[5]  & n29136;
  assign n29138 =  a[5]  & ~n29136;
  assign n29139 = ~n29135 & ~n29138;
  assign n29140 = ~n29137 & n29139;
  assign n29141 = ~n29135 & ~n29140;
  assign n29142 = ~n29138 & ~n29140;
  assign n29143 = ~n29137 & n29142;
  assign n29144 = ~n29141 & ~n29143;
  assign n29145 = ~n28925 & n29144;
  assign n29146 = n28925 & ~n29144;
  assign n29147 = ~n29145 & ~n29146;
  assign n29148 = n75 & n23368;
  assign n29149 = n3020 & n22359;
  assign n29150 = n3023 & n22365;
  assign n29151 = n3028 & n22362;
  assign n29152 = ~n29150 & ~n29151;
  assign n29153 = ~n29149 & n29152;
  assign n29154 = ~n29148 & n29153;
  assign n29155 = ~n29147 & ~n29154;
  assign n29156 = n29147 & n29154;
  assign n29157 = ~n29155 & ~n29156;
  assign n29158 = n29117 & ~n29157;
  assign n29159 = ~n29117 & n29157;
  assign n29160 = ~n29158 & ~n29159;
  assign n29161 = n3457 & n22350;
  assign n29162 = n3542 & n22356;
  assign n29163 = n3606 & n22353;
  assign n29164 = ~n29162 & ~n29163;
  assign n29165 = ~n29161 & n29164;
  assign n29166 = n3368 & n23672;
  assign n29167 = n29165 & ~n29166;
  assign n29168 =  a[29]  & ~n29167;
  assign n29169 =  a[29]  & ~n29168;
  assign n29170 = ~n29167 & ~n29168;
  assign n29171 = ~n29169 & ~n29170;
  assign n29172 = n29160 & ~n29171;
  assign n29173 = n29160 & ~n29172;
  assign n29174 = ~n29171 & ~n29172;
  assign n29175 = ~n29173 & ~n29174;
  assign n29176 = n3884 & n22341;
  assign n29177 = n3967 & n22347;
  assign n29178 = n4046 & n22344;
  assign n29179 = ~n29177 & ~n29178;
  assign n29180 = ~n29176 & n29179;
  assign n29181 = n4050 & n24142;
  assign n29182 = n29180 & ~n29181;
  assign n29183 =  a[26]  & ~n29182;
  assign n29184 =  a[26]  & ~n29183;
  assign n29185 = ~n29182 & ~n29183;
  assign n29186 = ~n29184 & ~n29185;
  assign n29187 = ~n29175 & ~n29186;
  assign n29188 = ~n29175 & ~n29187;
  assign n29189 = ~n29186 & ~n29187;
  assign n29190 = ~n29188 & ~n29189;
  assign n29191 = ~n28954 & ~n28969;
  assign n29192 = n29190 & n29191;
  assign n29193 = ~n29190 & ~n29191;
  assign n29194 = ~n29192 & ~n29193;
  assign n29195 = n4694 & n22332;
  assign n29196 = n4533 & n22338;
  assign n29197 = n4604 & n22335;
  assign n29198 = ~n29196 & ~n29197;
  assign n29199 = ~n29195 & n29198;
  assign n29200 = n4536 & n22542;
  assign n29201 = n29199 & ~n29200;
  assign n29202 =  a[23]  & ~n29201;
  assign n29203 =  a[23]  & ~n29202;
  assign n29204 = ~n29201 & ~n29202;
  assign n29205 = ~n29203 & ~n29204;
  assign n29206 = n29194 & ~n29205;
  assign n29207 = n29194 & ~n29206;
  assign n29208 = ~n29205 & ~n29206;
  assign n29209 = ~n29207 & ~n29208;
  assign n29210 = ~n28975 & ~n28988;
  assign n29211 = n29209 & n29210;
  assign n29212 = ~n29209 & ~n29210;
  assign n29213 = ~n29211 & ~n29212;
  assign n29214 = n5496 & n22323;
  assign n29215 = n4935 & n22329;
  assign n29216 = n5407 & n22326;
  assign n29217 = ~n29215 & ~n29216;
  assign n29218 = ~n29214 & n29217;
  assign n29219 = n4938 & n24599;
  assign n29220 = n29218 & ~n29219;
  assign n29221 =  a[20]  & ~n29220;
  assign n29222 =  a[20]  & ~n29221;
  assign n29223 = ~n29220 & ~n29221;
  assign n29224 = ~n29222 & ~n29223;
  assign n29225 = n29213 & ~n29224;
  assign n29226 = n29213 & ~n29225;
  assign n29227 = ~n29224 & ~n29225;
  assign n29228 = ~n29226 & ~n29227;
  assign n29229 = ~n28994 & ~n29007;
  assign n29230 = n29228 & n29229;
  assign n29231 = ~n29228 & ~n29229;
  assign n29232 = ~n29230 & ~n29231;
  assign n29233 = n6233 & n22315;
  assign n29234 = n5663 & n22320;
  assign n29235 = n5939 & n22312;
  assign n29236 = ~n29234 & ~n29235;
  assign n29237 = ~n29233 & n29236;
  assign n29238 = n5666 & n25294;
  assign n29239 = n29237 & ~n29238;
  assign n29240 =  a[17]  & ~n29239;
  assign n29241 =  a[17]  & ~n29240;
  assign n29242 = ~n29239 & ~n29240;
  assign n29243 = ~n29241 & ~n29242;
  assign n29244 = n29232 & ~n29243;
  assign n29245 = n29232 & ~n29244;
  assign n29246 = ~n29243 & ~n29244;
  assign n29247 = ~n29245 & ~n29246;
  assign n29248 = ~n29013 & ~n29026;
  assign n29249 = n29247 & n29248;
  assign n29250 = ~n29247 & ~n29248;
  assign n29251 = ~n29249 & ~n29250;
  assign n29252 = ~n29032 & ~n29045;
  assign n29253 = n7101 & n26066;
  assign n29254 = n6402 & n22309;
  assign n29255 = n6951 & n26063;
  assign n29256 = ~n29254 & ~n29255;
  assign n29257 = ~n29253 & n29256;
  assign n29258 = n6397 & ~n26624;
  assign n29259 = n29257 & ~n29258;
  assign n29260 =  a[14]  & ~n29259;
  assign n29261 =  a[14]  & ~n29260;
  assign n29262 = ~n29259 & ~n29260;
  assign n29263 = ~n29261 & ~n29262;
  assign n29264 = ~n29252 & ~n29263;
  assign n29265 = ~n29252 & ~n29264;
  assign n29266 = ~n29263 & ~n29264;
  assign n29267 = ~n29265 & ~n29266;
  assign n29268 = ~n29251 & n29267;
  assign n29269 = n29251 & ~n29267;
  assign n29270 = ~n29268 & ~n29269;
  assign n29271 = n7983 & n27173;
  assign n29272 = n7291 & n26060;
  assign n29273 = n7632 & n26890;
  assign n29274 = ~n29272 & ~n29273;
  assign n29275 = ~n29271 & n29274;
  assign n29276 = n7294 & n27185;
  assign n29277 = n29275 & ~n29276;
  assign n29278 =  a[11]  & ~n29277;
  assign n29279 =  a[11]  & ~n29278;
  assign n29280 = ~n29277 & ~n29278;
  assign n29281 = ~n29279 & ~n29280;
  assign n29282 = n29270 & ~n29281;
  assign n29283 = n29270 & ~n29282;
  assign n29284 = ~n29281 & ~n29282;
  assign n29285 = ~n29283 & ~n29284;
  assign n29286 = ~n29051 & ~n29064;
  assign n29287 = n29285 & n29286;
  assign n29288 = ~n29285 & ~n29286;
  assign n29289 = ~n29287 & ~n29288;
  assign n29290 = ~n29070 & ~n29083;
  assign n29291 = n9331 & n27964;
  assign n29292 = n8418 & n27442;
  assign n29293 = n8860 & n27698;
  assign n29294 = ~n29292 & ~n29293;
  assign n29295 = ~n29291 & n29294;
  assign n29296 = n8421 & n27976;
  assign n29297 = n29295 & ~n29296;
  assign n29298 =  a[8]  & ~n29297;
  assign n29299 =  a[8]  & ~n29298;
  assign n29300 = ~n29297 & ~n29298;
  assign n29301 = ~n29299 & ~n29300;
  assign n29302 = ~n29290 & ~n29301;
  assign n29303 = ~n29290 & ~n29302;
  assign n29304 = ~n29301 & ~n29302;
  assign n29305 = ~n29303 & ~n29304;
  assign n29306 = ~n29289 & n29305;
  assign n29307 = n29289 & ~n29305;
  assign n29308 = ~n29306 & ~n29307;
  assign n29309 = ~n29116 & n29308;
  assign n29310 = n29116 & ~n29308;
  assign n29311 = ~n29309 & ~n29310;
  assign n29312 = ~n29115 & n29311;
  assign n29313 = n29115 & ~n29311;
  assign n29314 = ~n29312 & ~n29313;
  assign n29315 = ~n29112 & ~n29314;
  assign n29316 = n29112 & n29314;
  assign  result[10]  = ~n29315 & ~n29316;
  assign n29318 = ~n29159 & ~n29172;
  assign n29319 = n75 & ~n23345;
  assign n29320 = n3020 & n22356;
  assign n29321 = n3023 & n22362;
  assign n29322 = n3028 & n22359;
  assign n29323 = ~n29321 & ~n29322;
  assign n29324 = ~n29320 & n29323;
  assign n29325 = ~n29319 & n29324;
  assign n29326 = n1324 & n6056;
  assign n29327 = n1206 & n29326;
  assign n29328 = n1346 & n29327;
  assign n29329 = n6705 & n29328;
  assign n29330 = n654 & n29329;
  assign n29331 = n3470 & n29330;
  assign n29332 = n869 & n29331;
  assign n29333 = n1141 & n29332;
  assign n29334 = ~n229 & n29333;
  assign n29335 = ~n121 & n29334;
  assign n29336 = ~n248 & n29335;
  assign n29337 = ~n206 & n29336;
  assign n29338 = n1732 & n2263;
  assign n29339 = n3160 & n29338;
  assign n29340 = n6771 & n29339;
  assign n29341 = n29337 & n29340;
  assign n29342 = n1378 & n29341;
  assign n29343 = n2678 & n29342;
  assign n29344 = n600 & n29343;
  assign n29345 = n488 & n29344;
  assign n29346 = n1009 & n29345;
  assign n29347 = n1825 & n29346;
  assign n29348 = n1522 & n29347;
  assign n29349 = ~n1011 & n29348;
  assign n29350 = ~n1246 & n29349;
  assign n29351 = ~n275 & n29350;
  assign n29352 = ~n357 & n29351;
  assign n29353 = ~n165 & n29352;
  assign n29354 = ~n493 & n29353;
  assign n29355 = ~n655 & n29354;
  assign n29356 = n28496 & ~n29132;
  assign n29357 = ~n29140 & ~n29356;
  assign n29358 = n29355 & ~n29357;
  assign n29359 = ~n29355 & n29357;
  assign n29360 = ~n29358 & ~n29359;
  assign n29361 = ~n29325 & n29360;
  assign n29362 = ~n29325 & ~n29361;
  assign n29363 = n29360 & ~n29361;
  assign n29364 = ~n29362 & ~n29363;
  assign n29365 = ~n28925 & ~n29144;
  assign n29366 = ~n29155 & ~n29365;
  assign n29367 = n29364 & n29366;
  assign n29368 = ~n29364 & ~n29366;
  assign n29369 = ~n29367 & ~n29368;
  assign n29370 = n3457 & n22347;
  assign n29371 = n3542 & n22353;
  assign n29372 = n3606 & n22350;
  assign n29373 = ~n29371 & ~n29372;
  assign n29374 = ~n29370 & n29373;
  assign n29375 = ~n3368 & n29374;
  assign n29376 = n23659 & n29374;
  assign n29377 = ~n29375 & ~n29376;
  assign n29378 =  a[29]  & ~n29377;
  assign n29379 = ~ a[29]  & n29377;
  assign n29380 = ~n29378 & ~n29379;
  assign n29381 = n29369 & ~n29380;
  assign n29382 = ~n29369 & n29380;
  assign n29383 = ~n29381 & ~n29382;
  assign n29384 = ~n29318 & n29383;
  assign n29385 = n29318 & ~n29383;
  assign n29386 = ~n29384 & ~n29385;
  assign n29387 = n3884 & n22338;
  assign n29388 = n3967 & n22344;
  assign n29389 = n4046 & n22341;
  assign n29390 = ~n29388 & ~n29389;
  assign n29391 = ~n29387 & n29390;
  assign n29392 = n4050 & ~n24188;
  assign n29393 = n29391 & ~n29392;
  assign n29394 =  a[26]  & ~n29393;
  assign n29395 =  a[26]  & ~n29394;
  assign n29396 = ~n29393 & ~n29394;
  assign n29397 = ~n29395 & ~n29396;
  assign n29398 = n29386 & ~n29397;
  assign n29399 = n29386 & ~n29398;
  assign n29400 = ~n29397 & ~n29398;
  assign n29401 = ~n29399 & ~n29400;
  assign n29402 = ~n29187 & ~n29193;
  assign n29403 = n29401 & n29402;
  assign n29404 = ~n29401 & ~n29402;
  assign n29405 = ~n29403 & ~n29404;
  assign n29406 = n4694 & n22329;
  assign n29407 = n4533 & n22335;
  assign n29408 = n4604 & n22332;
  assign n29409 = ~n29407 & ~n29408;
  assign n29410 = ~n29406 & n29409;
  assign n29411 = n4536 & ~n24633;
  assign n29412 = n29410 & ~n29411;
  assign n29413 =  a[23]  & ~n29412;
  assign n29414 =  a[23]  & ~n29413;
  assign n29415 = ~n29412 & ~n29413;
  assign n29416 = ~n29414 & ~n29415;
  assign n29417 = n29405 & ~n29416;
  assign n29418 = n29405 & ~n29417;
  assign n29419 = ~n29416 & ~n29417;
  assign n29420 = ~n29418 & ~n29419;
  assign n29421 = ~n29206 & ~n29212;
  assign n29422 = n29420 & n29421;
  assign n29423 = ~n29420 & ~n29421;
  assign n29424 = ~n29422 & ~n29423;
  assign n29425 = n5496 & n22320;
  assign n29426 = n4935 & n22326;
  assign n29427 = n5407 & n22323;
  assign n29428 = ~n29426 & ~n29427;
  assign n29429 = ~n29425 & n29428;
  assign n29430 = n4938 & ~n25270;
  assign n29431 = n29429 & ~n29430;
  assign n29432 =  a[20]  & ~n29431;
  assign n29433 =  a[20]  & ~n29432;
  assign n29434 = ~n29431 & ~n29432;
  assign n29435 = ~n29433 & ~n29434;
  assign n29436 = n29424 & ~n29435;
  assign n29437 = n29424 & ~n29436;
  assign n29438 = ~n29435 & ~n29436;
  assign n29439 = ~n29437 & ~n29438;
  assign n29440 = ~n29225 & ~n29231;
  assign n29441 = n29439 & n29440;
  assign n29442 = ~n29439 & ~n29440;
  assign n29443 = ~n29441 & ~n29442;
  assign n29444 = n6233 & n22309;
  assign n29445 = n5663 & n22312;
  assign n29446 = n5939 & n22315;
  assign n29447 = ~n29445 & ~n29446;
  assign n29448 = ~n29444 & n29447;
  assign n29449 = n5666 & ~n22529;
  assign n29450 = n29448 & ~n29449;
  assign n29451 =  a[17]  & ~n29450;
  assign n29452 =  a[17]  & ~n29451;
  assign n29453 = ~n29450 & ~n29451;
  assign n29454 = ~n29452 & ~n29453;
  assign n29455 = n29443 & ~n29454;
  assign n29456 = n29443 & ~n29455;
  assign n29457 = ~n29454 & ~n29455;
  assign n29458 = ~n29456 & ~n29457;
  assign n29459 = ~n29244 & ~n29250;
  assign n29460 = n29458 & n29459;
  assign n29461 = ~n29458 & ~n29459;
  assign n29462 = ~n29460 & ~n29461;
  assign n29463 = n7101 & n26060;
  assign n29464 = n6402 & n26063;
  assign n29465 = n6951 & n26066;
  assign n29466 = ~n29464 & ~n29465;
  assign n29467 = ~n29463 & n29466;
  assign n29468 = n6397 & ~n26088;
  assign n29469 = n29467 & ~n29468;
  assign n29470 =  a[14]  & ~n29469;
  assign n29471 =  a[14]  & ~n29470;
  assign n29472 = ~n29469 & ~n29470;
  assign n29473 = ~n29471 & ~n29472;
  assign n29474 = n29462 & ~n29473;
  assign n29475 = n29462 & ~n29474;
  assign n29476 = ~n29473 & ~n29474;
  assign n29477 = ~n29475 & ~n29476;
  assign n29478 = ~n29264 & ~n29269;
  assign n29479 = ~n29477 & ~n29478;
  assign n29480 = ~n29477 & ~n29479;
  assign n29481 = ~n29478 & ~n29479;
  assign n29482 = ~n29480 & ~n29481;
  assign n29483 = n7983 & n27442;
  assign n29484 = n7291 & n26890;
  assign n29485 = n7632 & n27173;
  assign n29486 = ~n29484 & ~n29485;
  assign n29487 = ~n29483 & n29486;
  assign n29488 = n7294 & n27455;
  assign n29489 = n29487 & ~n29488;
  assign n29490 =  a[11]  & ~n29489;
  assign n29491 =  a[11]  & ~n29490;
  assign n29492 = ~n29489 & ~n29490;
  assign n29493 = ~n29491 & ~n29492;
  assign n29494 = ~n29482 & ~n29493;
  assign n29495 = ~n29482 & ~n29494;
  assign n29496 = ~n29493 & ~n29494;
  assign n29497 = ~n29495 & ~n29496;
  assign n29498 = ~n29282 & ~n29288;
  assign n29499 = n29497 & n29498;
  assign n29500 = ~n29497 & ~n29498;
  assign n29501 = ~n29499 & ~n29500;
  assign n29502 = n9331 & ~n28208;
  assign n29503 = n8418 & n27698;
  assign n29504 = n8860 & n27964;
  assign n29505 = ~n29503 & ~n29504;
  assign n29506 = ~n29502 & n29505;
  assign n29507 = n8421 & ~n28223;
  assign n29508 = n29506 & ~n29507;
  assign n29509 =  a[8]  & ~n29508;
  assign n29510 =  a[8]  & ~n29509;
  assign n29511 = ~n29508 & ~n29509;
  assign n29512 = ~n29510 & ~n29511;
  assign n29513 = n29501 & ~n29512;
  assign n29514 = n29501 & ~n29513;
  assign n29515 = ~n29512 & ~n29513;
  assign n29516 = ~n29514 & ~n29515;
  assign n29517 = ~n29302 & ~n29307;
  assign n29518 = ~n29516 & ~n29517;
  assign n29519 = ~n29516 & ~n29518;
  assign n29520 = ~n29517 & ~n29518;
  assign n29521 = ~n29519 & ~n29520;
  assign n29522 = ~n29309 & ~n29312;
  assign n29523 = n29521 & n29522;
  assign n29524 = ~n29521 & ~n29522;
  assign n29525 = ~n29523 & ~n29524;
  assign n29526 = ~n29316 & n29525;
  assign n29527 = n29316 & ~n29525;
  assign  result[11]  = n29526 | n29527;
  assign n29529 = n29316 & n29525;
  assign n29530 = ~n29358 & ~n29361;
  assign n29531 = ~n175 & ~n255;
  assign n29532 = ~n299 & n29531;
  assign n29533 = ~n305 & n29532;
  assign n29534 = ~n492 & n29533;
  assign n29535 = ~n165 & n29534;
  assign n29536 = ~n592 & n29535;
  assign n29537 = ~n672 & n29536;
  assign n29538 = ~n270 & n29537;
  assign n29539 = n2442 & n12712;
  assign n29540 = n940 & n29539;
  assign n29541 = n4295 & n29540;
  assign n29542 = n2406 & n29541;
  assign n29543 = n1046 & n29542;
  assign n29544 = n2417 & n29543;
  assign n29545 = n885 & n29544;
  assign n29546 = ~n289 & n29545;
  assign n29547 = ~n155 & n29546;
  assign n29548 = ~n164 & n29547;
  assign n29549 = ~n191 & n29548;
  assign n29550 = ~n245 & n29549;
  assign n29551 = n12911 & n13808;
  assign n29552 = n6548 & n29551;
  assign n29553 = n29550 & n29552;
  assign n29554 = n29538 & n29553;
  assign n29555 = n3065 & n29554;
  assign n29556 = n12396 & n29555;
  assign n29557 = ~n194 & n29556;
  assign n29558 = ~n254 & n29557;
  assign n29559 = ~n435 & n29558;
  assign n29560 = ~n243 & n29559;
  assign n29561 = ~n466 & n29560;
  assign n29562 = ~n537 & n29561;
  assign n29563 = ~n332 & n29562;
  assign n29564 = ~n325 & n29563;
  assign n29565 = ~n29355 & n29564;
  assign n29566 = n29355 & ~n29564;
  assign n29567 = ~n29530 & ~n29566;
  assign n29568 = ~n29565 & n29567;
  assign n29569 = ~n29530 & ~n29568;
  assign n29570 = ~n29566 & ~n29568;
  assign n29571 = ~n29565 & n29570;
  assign n29572 = ~n29569 & ~n29571;
  assign n29573 = n75 & ~n22556;
  assign n29574 = n3020 & n22353;
  assign n29575 = n3023 & n22359;
  assign n29576 = n3028 & n22356;
  assign n29577 = ~n29575 & ~n29576;
  assign n29578 = ~n29574 & n29577;
  assign n29579 = ~n29573 & n29578;
  assign n29580 = ~n29572 & ~n29579;
  assign n29581 = ~n29572 & ~n29580;
  assign n29582 = ~n29579 & ~n29580;
  assign n29583 = ~n29581 & ~n29582;
  assign n29584 = ~n29368 & ~n29381;
  assign n29585 = n29583 & n29584;
  assign n29586 = ~n29583 & ~n29584;
  assign n29587 = ~n29585 & ~n29586;
  assign n29588 = n3457 & n22344;
  assign n29589 = n3542 & n22350;
  assign n29590 = n3606 & n22347;
  assign n29591 = ~n29589 & ~n29590;
  assign n29592 = ~n29588 & n29591;
  assign n29593 = n3368 & ~n23642;
  assign n29594 = n29592 & ~n29593;
  assign n29595 =  a[29]  & ~n29594;
  assign n29596 =  a[29]  & ~n29595;
  assign n29597 = ~n29594 & ~n29595;
  assign n29598 = ~n29596 & ~n29597;
  assign n29599 = n29587 & ~n29598;
  assign n29600 = n29587 & ~n29599;
  assign n29601 = ~n29598 & ~n29599;
  assign n29602 = ~n29600 & ~n29601;
  assign n29603 = n3884 & n22335;
  assign n29604 = n3967 & n22341;
  assign n29605 = n4046 & n22338;
  assign n29606 = ~n29604 & ~n29605;
  assign n29607 = ~n29603 & n29606;
  assign n29608 = n4050 & ~n24167;
  assign n29609 = n29607 & ~n29608;
  assign n29610 =  a[26]  & ~n29609;
  assign n29611 =  a[26]  & ~n29610;
  assign n29612 = ~n29609 & ~n29610;
  assign n29613 = ~n29611 & ~n29612;
  assign n29614 = ~n29602 & ~n29613;
  assign n29615 = ~n29602 & ~n29614;
  assign n29616 = ~n29613 & ~n29614;
  assign n29617 = ~n29615 & ~n29616;
  assign n29618 = ~n29384 & ~n29398;
  assign n29619 = n29617 & n29618;
  assign n29620 = ~n29617 & ~n29618;
  assign n29621 = ~n29619 & ~n29620;
  assign n29622 = n4694 & n22326;
  assign n29623 = n4533 & n22332;
  assign n29624 = n4604 & n22329;
  assign n29625 = ~n29623 & ~n29624;
  assign n29626 = ~n29622 & n29625;
  assign n29627 = n4536 & ~n24616;
  assign n29628 = n29626 & ~n29627;
  assign n29629 =  a[23]  & ~n29628;
  assign n29630 =  a[23]  & ~n29629;
  assign n29631 = ~n29628 & ~n29629;
  assign n29632 = ~n29630 & ~n29631;
  assign n29633 = n29621 & ~n29632;
  assign n29634 = n29621 & ~n29633;
  assign n29635 = ~n29632 & ~n29633;
  assign n29636 = ~n29634 & ~n29635;
  assign n29637 = ~n29404 & ~n29417;
  assign n29638 = n29636 & n29637;
  assign n29639 = ~n29636 & ~n29637;
  assign n29640 = ~n29638 & ~n29639;
  assign n29641 = n5496 & n22312;
  assign n29642 = n4935 & n22323;
  assign n29643 = n5407 & n22320;
  assign n29644 = ~n29642 & ~n29643;
  assign n29645 = ~n29641 & n29644;
  assign n29646 = n4938 & ~n25315;
  assign n29647 = n29645 & ~n29646;
  assign n29648 =  a[20]  & ~n29647;
  assign n29649 =  a[20]  & ~n29648;
  assign n29650 = ~n29647 & ~n29648;
  assign n29651 = ~n29649 & ~n29650;
  assign n29652 = n29640 & ~n29651;
  assign n29653 = n29640 & ~n29652;
  assign n29654 = ~n29651 & ~n29652;
  assign n29655 = ~n29653 & ~n29654;
  assign n29656 = ~n29423 & ~n29436;
  assign n29657 = n29655 & n29656;
  assign n29658 = ~n29655 & ~n29656;
  assign n29659 = ~n29657 & ~n29658;
  assign n29660 = n6233 & n26063;
  assign n29661 = n5663 & n22315;
  assign n29662 = n5939 & n22309;
  assign n29663 = ~n29661 & ~n29662;
  assign n29664 = ~n29660 & n29663;
  assign n29665 = n5666 & ~n26604;
  assign n29666 = n29664 & ~n29665;
  assign n29667 =  a[17]  & ~n29666;
  assign n29668 =  a[17]  & ~n29667;
  assign n29669 = ~n29666 & ~n29667;
  assign n29670 = ~n29668 & ~n29669;
  assign n29671 = n29659 & ~n29670;
  assign n29672 = n29659 & ~n29671;
  assign n29673 = ~n29670 & ~n29671;
  assign n29674 = ~n29672 & ~n29673;
  assign n29675 = ~n29442 & ~n29455;
  assign n29676 = n29674 & n29675;
  assign n29677 = ~n29674 & ~n29675;
  assign n29678 = ~n29676 & ~n29677;
  assign n29679 = n7101 & n26890;
  assign n29680 = n6402 & n26066;
  assign n29681 = n6951 & n26060;
  assign n29682 = ~n29680 & ~n29681;
  assign n29683 = ~n29679 & n29682;
  assign n29684 = n6397 & ~n26904;
  assign n29685 = n29683 & ~n29684;
  assign n29686 =  a[14]  & ~n29685;
  assign n29687 =  a[14]  & ~n29686;
  assign n29688 = ~n29685 & ~n29686;
  assign n29689 = ~n29687 & ~n29688;
  assign n29690 = n29678 & ~n29689;
  assign n29691 = n29678 & ~n29690;
  assign n29692 = ~n29689 & ~n29690;
  assign n29693 = ~n29691 & ~n29692;
  assign n29694 = ~n29461 & ~n29474;
  assign n29695 = n29693 & n29694;
  assign n29696 = ~n29693 & ~n29694;
  assign n29697 = ~n29695 & ~n29696;
  assign n29698 = n7983 & n27698;
  assign n29699 = n7291 & n27173;
  assign n29700 = n7632 & n27442;
  assign n29701 = ~n29699 & ~n29700;
  assign n29702 = ~n29698 & n29701;
  assign n29703 = n7294 & ~n27713;
  assign n29704 = n29702 & ~n29703;
  assign n29705 =  a[11]  & ~n29704;
  assign n29706 =  a[11]  & ~n29705;
  assign n29707 = ~n29704 & ~n29705;
  assign n29708 = ~n29706 & ~n29707;
  assign n29709 = n29697 & ~n29708;
  assign n29710 = n29697 & ~n29709;
  assign n29711 = ~n29708 & ~n29709;
  assign n29712 = ~n29710 & ~n29711;
  assign n29713 = ~n29479 & ~n29494;
  assign n29714 = ~n14590 & ~n28208;
  assign n29715 = n8418 & n27964;
  assign n29716 = ~n29714 & ~n29715;
  assign n29717 = ~n8421 & n29716;
  assign n29718 = n28221 & n29716;
  assign n29719 = ~n29717 & ~n29718;
  assign n29720 =  a[8]  & ~n29719;
  assign n29721 = ~ a[8]  & n29719;
  assign n29722 = ~n29720 & ~n29721;
  assign n29723 = ~n29713 & ~n29722;
  assign n29724 = n29713 & n29722;
  assign n29725 = ~n29723 & ~n29724;
  assign n29726 = ~n29712 & n29725;
  assign n29727 = ~n29712 & ~n29726;
  assign n29728 = n29725 & ~n29726;
  assign n29729 = ~n29727 & ~n29728;
  assign n29730 = ~n29500 & ~n29513;
  assign n29731 = n29729 & n29730;
  assign n29732 = ~n29729 & ~n29730;
  assign n29733 = ~n29731 & ~n29732;
  assign n29734 = ~n29518 & ~n29524;
  assign n29735 = ~n29733 & n29734;
  assign n29736 = n29733 & ~n29734;
  assign n29737 = ~n29735 & ~n29736;
  assign n29738 = n29529 & n29737;
  assign n29739 = ~n29529 & ~n29737;
  assign  result[12]  = ~n29738 & ~n29739;
  assign n29741 = ~n29732 & ~n29736;
  assign n29742 = ~n29723 & ~n29726;
  assign n29743 = n75 & n23672;
  assign n29744 = n3020 & n22350;
  assign n29745 = n3023 & n22356;
  assign n29746 = n3028 & n22353;
  assign n29747 = ~n29745 & ~n29746;
  assign n29748 = ~n29744 & n29747;
  assign n29749 = ~n29743 & n29748;
  assign n29750 = ~n14592 & ~n28208;
  assign n29751 =  a[8]  & ~n29750;
  assign n29752 = ~ a[8]  & n29750;
  assign n29753 = ~n29751 & ~n29752;
  assign n29754 = n960 & n3474;
  assign n29755 = n1422 & n29754;
  assign n29756 = n300 & n29755;
  assign n29757 = n13773 & n29756;
  assign n29758 = n2006 & n29757;
  assign n29759 = n1575 & n29758;
  assign n29760 = n2697 & n29759;
  assign n29761 = n235 & n29760;
  assign n29762 = n2958 & n29761;
  assign n29763 = n2484 & n29762;
  assign n29764 = n2170 & n29763;
  assign n29765 = n156 & n29764;
  assign n29766 = ~n713 & n29765;
  assign n29767 = ~n368 & n29766;
  assign n29768 = n29355 & n29767;
  assign n29769 = ~n29355 & ~n29767;
  assign n29770 = ~n29768 & ~n29769;
  assign n29771 = n29753 & n29770;
  assign n29772 = ~n29753 & ~n29770;
  assign n29773 = ~n29771 & ~n29772;
  assign n29774 = ~n29570 & n29773;
  assign n29775 = n29570 & ~n29773;
  assign n29776 = ~n29774 & ~n29775;
  assign n29777 = ~n29749 & n29776;
  assign n29778 = n29776 & ~n29777;
  assign n29779 = ~n29749 & ~n29777;
  assign n29780 = ~n29778 & ~n29779;
  assign n29781 = n3457 & n22341;
  assign n29782 = n3542 & n22347;
  assign n29783 = n3606 & n22344;
  assign n29784 = ~n29782 & ~n29783;
  assign n29785 = ~n29781 & n29784;
  assign n29786 = n3368 & n24142;
  assign n29787 = n29785 & ~n29786;
  assign n29788 =  a[29]  & ~n29787;
  assign n29789 =  a[29]  & ~n29788;
  assign n29790 = ~n29787 & ~n29788;
  assign n29791 = ~n29789 & ~n29790;
  assign n29792 = ~n29780 & ~n29791;
  assign n29793 = ~n29780 & ~n29792;
  assign n29794 = ~n29791 & ~n29792;
  assign n29795 = ~n29793 & ~n29794;
  assign n29796 = ~n29580 & ~n29586;
  assign n29797 = n29795 & n29796;
  assign n29798 = ~n29795 & ~n29796;
  assign n29799 = ~n29797 & ~n29798;
  assign n29800 = n3884 & n22332;
  assign n29801 = n3967 & n22338;
  assign n29802 = n4046 & n22335;
  assign n29803 = ~n29801 & ~n29802;
  assign n29804 = ~n29800 & n29803;
  assign n29805 = n4050 & n22542;
  assign n29806 = n29804 & ~n29805;
  assign n29807 =  a[26]  & ~n29806;
  assign n29808 =  a[26]  & ~n29807;
  assign n29809 = ~n29806 & ~n29807;
  assign n29810 = ~n29808 & ~n29809;
  assign n29811 = n29799 & ~n29810;
  assign n29812 = n29799 & ~n29811;
  assign n29813 = ~n29810 & ~n29811;
  assign n29814 = ~n29812 & ~n29813;
  assign n29815 = ~n29599 & ~n29614;
  assign n29816 = n29814 & n29815;
  assign n29817 = ~n29814 & ~n29815;
  assign n29818 = ~n29816 & ~n29817;
  assign n29819 = n4694 & n22323;
  assign n29820 = n4533 & n22329;
  assign n29821 = n4604 & n22326;
  assign n29822 = ~n29820 & ~n29821;
  assign n29823 = ~n29819 & n29822;
  assign n29824 = n4536 & n24599;
  assign n29825 = n29823 & ~n29824;
  assign n29826 =  a[23]  & ~n29825;
  assign n29827 =  a[23]  & ~n29826;
  assign n29828 = ~n29825 & ~n29826;
  assign n29829 = ~n29827 & ~n29828;
  assign n29830 = n29818 & ~n29829;
  assign n29831 = n29818 & ~n29830;
  assign n29832 = ~n29829 & ~n29830;
  assign n29833 = ~n29831 & ~n29832;
  assign n29834 = ~n29620 & ~n29633;
  assign n29835 = n29833 & n29834;
  assign n29836 = ~n29833 & ~n29834;
  assign n29837 = ~n29835 & ~n29836;
  assign n29838 = n5496 & n22315;
  assign n29839 = n4935 & n22320;
  assign n29840 = n5407 & n22312;
  assign n29841 = ~n29839 & ~n29840;
  assign n29842 = ~n29838 & n29841;
  assign n29843 = n4938 & n25294;
  assign n29844 = n29842 & ~n29843;
  assign n29845 =  a[20]  & ~n29844;
  assign n29846 =  a[20]  & ~n29845;
  assign n29847 = ~n29844 & ~n29845;
  assign n29848 = ~n29846 & ~n29847;
  assign n29849 = n29837 & ~n29848;
  assign n29850 = n29837 & ~n29849;
  assign n29851 = ~n29848 & ~n29849;
  assign n29852 = ~n29850 & ~n29851;
  assign n29853 = ~n29639 & ~n29652;
  assign n29854 = n29852 & n29853;
  assign n29855 = ~n29852 & ~n29853;
  assign n29856 = ~n29854 & ~n29855;
  assign n29857 = ~n29658 & ~n29671;
  assign n29858 = n6233 & n26066;
  assign n29859 = n5663 & n22309;
  assign n29860 = n5939 & n26063;
  assign n29861 = ~n29859 & ~n29860;
  assign n29862 = ~n29858 & n29861;
  assign n29863 = n5666 & ~n26624;
  assign n29864 = n29862 & ~n29863;
  assign n29865 =  a[17]  & ~n29864;
  assign n29866 =  a[17]  & ~n29865;
  assign n29867 = ~n29864 & ~n29865;
  assign n29868 = ~n29866 & ~n29867;
  assign n29869 = ~n29857 & ~n29868;
  assign n29870 = ~n29857 & ~n29869;
  assign n29871 = ~n29868 & ~n29869;
  assign n29872 = ~n29870 & ~n29871;
  assign n29873 = ~n29856 & n29872;
  assign n29874 = n29856 & ~n29872;
  assign n29875 = ~n29873 & ~n29874;
  assign n29876 = n7101 & n27173;
  assign n29877 = n6402 & n26060;
  assign n29878 = n6951 & n26890;
  assign n29879 = ~n29877 & ~n29878;
  assign n29880 = ~n29876 & n29879;
  assign n29881 = n6397 & n27185;
  assign n29882 = n29880 & ~n29881;
  assign n29883 =  a[14]  & ~n29882;
  assign n29884 =  a[14]  & ~n29883;
  assign n29885 = ~n29882 & ~n29883;
  assign n29886 = ~n29884 & ~n29885;
  assign n29887 = n29875 & ~n29886;
  assign n29888 = n29875 & ~n29887;
  assign n29889 = ~n29886 & ~n29887;
  assign n29890 = ~n29888 & ~n29889;
  assign n29891 = ~n29677 & ~n29690;
  assign n29892 = n29890 & n29891;
  assign n29893 = ~n29890 & ~n29891;
  assign n29894 = ~n29892 & ~n29893;
  assign n29895 = ~n29696 & ~n29709;
  assign n29896 = n7983 & n27964;
  assign n29897 = n7291 & n27442;
  assign n29898 = n7632 & n27698;
  assign n29899 = ~n29897 & ~n29898;
  assign n29900 = ~n29896 & n29899;
  assign n29901 = n7294 & n27976;
  assign n29902 = n29900 & ~n29901;
  assign n29903 =  a[11]  & ~n29902;
  assign n29904 =  a[11]  & ~n29903;
  assign n29905 = ~n29902 & ~n29903;
  assign n29906 = ~n29904 & ~n29905;
  assign n29907 = ~n29895 & ~n29906;
  assign n29908 = ~n29895 & ~n29907;
  assign n29909 = ~n29906 & ~n29907;
  assign n29910 = ~n29908 & ~n29909;
  assign n29911 = ~n29894 & n29910;
  assign n29912 = n29894 & ~n29910;
  assign n29913 = ~n29911 & ~n29912;
  assign n29914 = ~n29742 & n29913;
  assign n29915 = n29742 & ~n29913;
  assign n29916 = ~n29914 & ~n29915;
  assign n29917 = ~n29741 & n29916;
  assign n29918 = n29741 & ~n29916;
  assign n29919 = ~n29917 & ~n29918;
  assign n29920 = ~n29738 & ~n29919;
  assign n29921 = n29738 & n29919;
  assign  result[13]  = ~n29920 & ~n29921;
  assign n29923 = ~n29792 & ~n29798;
  assign n29924 = n75 & ~n23659;
  assign n29925 = n3020 & n22347;
  assign n29926 = n3023 & n22353;
  assign n29927 = n3028 & n22350;
  assign n29928 = ~n29926 & ~n29927;
  assign n29929 = ~n29925 & n29928;
  assign n29930 = ~n29924 & n29929;
  assign n29931 = ~n29769 & ~n29771;
  assign n29932 = n962 & n1490;
  assign n29933 = n15854 & n29932;
  assign n29934 = n14407 & n29933;
  assign n29935 = n4767 & n29934;
  assign n29936 = n4786 & n29935;
  assign n29937 = n1719 & n29936;
  assign n29938 = n3559 & n29937;
  assign n29939 = n2635 & n29938;
  assign n29940 = ~n242 & n29939;
  assign n29941 = ~n150 & n29940;
  assign n29942 = ~n357 & n29941;
  assign n29943 = ~n286 & n29942;
  assign n29944 = ~n980 & n29943;
  assign n29945 = ~n1010 & n29944;
  assign n29946 = ~n270 & n29945;
  assign n29947 = ~n29931 & n29946;
  assign n29948 = n29931 & ~n29946;
  assign n29949 = ~n29947 & ~n29948;
  assign n29950 = ~n29930 & n29949;
  assign n29951 = ~n29930 & ~n29950;
  assign n29952 = n29949 & ~n29950;
  assign n29953 = ~n29951 & ~n29952;
  assign n29954 = ~n29774 & ~n29777;
  assign n29955 = n29953 & n29954;
  assign n29956 = ~n29953 & ~n29954;
  assign n29957 = ~n29955 & ~n29956;
  assign n29958 = n3457 & n22338;
  assign n29959 = n3542 & n22344;
  assign n29960 = n3606 & n22341;
  assign n29961 = ~n29959 & ~n29960;
  assign n29962 = ~n29958 & n29961;
  assign n29963 = ~n3368 & n29962;
  assign n29964 = n24188 & n29962;
  assign n29965 = ~n29963 & ~n29964;
  assign n29966 =  a[29]  & ~n29965;
  assign n29967 = ~ a[29]  & n29965;
  assign n29968 = ~n29966 & ~n29967;
  assign n29969 = n29957 & ~n29968;
  assign n29970 = ~n29957 & n29968;
  assign n29971 = ~n29969 & ~n29970;
  assign n29972 = ~n29923 & n29971;
  assign n29973 = n29923 & ~n29971;
  assign n29974 = ~n29972 & ~n29973;
  assign n29975 = n3884 & n22329;
  assign n29976 = n3967 & n22335;
  assign n29977 = n4046 & n22332;
  assign n29978 = ~n29976 & ~n29977;
  assign n29979 = ~n29975 & n29978;
  assign n29980 = n4050 & ~n24633;
  assign n29981 = n29979 & ~n29980;
  assign n29982 =  a[26]  & ~n29981;
  assign n29983 =  a[26]  & ~n29982;
  assign n29984 = ~n29981 & ~n29982;
  assign n29985 = ~n29983 & ~n29984;
  assign n29986 = n29974 & ~n29985;
  assign n29987 = n29974 & ~n29986;
  assign n29988 = ~n29985 & ~n29986;
  assign n29989 = ~n29987 & ~n29988;
  assign n29990 = ~n29811 & ~n29817;
  assign n29991 = n29989 & n29990;
  assign n29992 = ~n29989 & ~n29990;
  assign n29993 = ~n29991 & ~n29992;
  assign n29994 = n4694 & n22320;
  assign n29995 = n4533 & n22326;
  assign n29996 = n4604 & n22323;
  assign n29997 = ~n29995 & ~n29996;
  assign n29998 = ~n29994 & n29997;
  assign n29999 = n4536 & ~n25270;
  assign n30000 = n29998 & ~n29999;
  assign n30001 =  a[23]  & ~n30000;
  assign n30002 =  a[23]  & ~n30001;
  assign n30003 = ~n30000 & ~n30001;
  assign n30004 = ~n30002 & ~n30003;
  assign n30005 = n29993 & ~n30004;
  assign n30006 = n29993 & ~n30005;
  assign n30007 = ~n30004 & ~n30005;
  assign n30008 = ~n30006 & ~n30007;
  assign n30009 = ~n29830 & ~n29836;
  assign n30010 = n30008 & n30009;
  assign n30011 = ~n30008 & ~n30009;
  assign n30012 = ~n30010 & ~n30011;
  assign n30013 = n5496 & n22309;
  assign n30014 = n4935 & n22312;
  assign n30015 = n5407 & n22315;
  assign n30016 = ~n30014 & ~n30015;
  assign n30017 = ~n30013 & n30016;
  assign n30018 = n4938 & ~n22529;
  assign n30019 = n30017 & ~n30018;
  assign n30020 =  a[20]  & ~n30019;
  assign n30021 =  a[20]  & ~n30020;
  assign n30022 = ~n30019 & ~n30020;
  assign n30023 = ~n30021 & ~n30022;
  assign n30024 = n30012 & ~n30023;
  assign n30025 = n30012 & ~n30024;
  assign n30026 = ~n30023 & ~n30024;
  assign n30027 = ~n30025 & ~n30026;
  assign n30028 = ~n29849 & ~n29855;
  assign n30029 = n30027 & n30028;
  assign n30030 = ~n30027 & ~n30028;
  assign n30031 = ~n30029 & ~n30030;
  assign n30032 = n6233 & n26060;
  assign n30033 = n5663 & n26063;
  assign n30034 = n5939 & n26066;
  assign n30035 = ~n30033 & ~n30034;
  assign n30036 = ~n30032 & n30035;
  assign n30037 = n5666 & ~n26088;
  assign n30038 = n30036 & ~n30037;
  assign n30039 =  a[17]  & ~n30038;
  assign n30040 =  a[17]  & ~n30039;
  assign n30041 = ~n30038 & ~n30039;
  assign n30042 = ~n30040 & ~n30041;
  assign n30043 = n30031 & ~n30042;
  assign n30044 = n30031 & ~n30043;
  assign n30045 = ~n30042 & ~n30043;
  assign n30046 = ~n30044 & ~n30045;
  assign n30047 = ~n29869 & ~n29874;
  assign n30048 = ~n30046 & ~n30047;
  assign n30049 = ~n30046 & ~n30048;
  assign n30050 = ~n30047 & ~n30048;
  assign n30051 = ~n30049 & ~n30050;
  assign n30052 = n7101 & n27442;
  assign n30053 = n6402 & n26890;
  assign n30054 = n6951 & n27173;
  assign n30055 = ~n30053 & ~n30054;
  assign n30056 = ~n30052 & n30055;
  assign n30057 = n6397 & n27455;
  assign n30058 = n30056 & ~n30057;
  assign n30059 =  a[14]  & ~n30058;
  assign n30060 =  a[14]  & ~n30059;
  assign n30061 = ~n30058 & ~n30059;
  assign n30062 = ~n30060 & ~n30061;
  assign n30063 = ~n30051 & ~n30062;
  assign n30064 = ~n30051 & ~n30063;
  assign n30065 = ~n30062 & ~n30063;
  assign n30066 = ~n30064 & ~n30065;
  assign n30067 = ~n29887 & ~n29893;
  assign n30068 = n30066 & n30067;
  assign n30069 = ~n30066 & ~n30067;
  assign n30070 = ~n30068 & ~n30069;
  assign n30071 = n7983 & ~n28208;
  assign n30072 = n7291 & n27698;
  assign n30073 = n7632 & n27964;
  assign n30074 = ~n30072 & ~n30073;
  assign n30075 = ~n30071 & n30074;
  assign n30076 = n7294 & ~n28223;
  assign n30077 = n30075 & ~n30076;
  assign n30078 =  a[11]  & ~n30077;
  assign n30079 =  a[11]  & ~n30078;
  assign n30080 = ~n30077 & ~n30078;
  assign n30081 = ~n30079 & ~n30080;
  assign n30082 = n30070 & ~n30081;
  assign n30083 = n30070 & ~n30082;
  assign n30084 = ~n30081 & ~n30082;
  assign n30085 = ~n30083 & ~n30084;
  assign n30086 = ~n29907 & ~n29912;
  assign n30087 = ~n30085 & ~n30086;
  assign n30088 = ~n30085 & ~n30087;
  assign n30089 = ~n30086 & ~n30087;
  assign n30090 = ~n30088 & ~n30089;
  assign n30091 = ~n29914 & ~n29917;
  assign n30092 = n30090 & n30091;
  assign n30093 = ~n30090 & ~n30091;
  assign n30094 = ~n30092 & ~n30093;
  assign n30095 = n29921 & ~n30094;
  assign n30096 = ~n29921 & n30094;
  assign  result[14]  = n30095 | n30096;
  assign n30098 = ~n29956 & ~n29969;
  assign n30099 = ~n29947 & ~n29950;
  assign n30100 = n2705 & n2811;
  assign n30101 = n2007 & n30100;
  assign n30102 = n1012 & n30101;
  assign n30103 = n877 & n30102;
  assign n30104 = n13768 & n30103;
  assign n30105 = n15312 & n30104;
  assign n30106 = n5286 & n30105;
  assign n30107 = n2651 & n30106;
  assign n30108 = n291 & n30107;
  assign n30109 = n1330 & n30108;
  assign n30110 = n29337 & n30109;
  assign n30111 = n731 & n30110;
  assign n30112 = n1247 & n30111;
  assign n30113 = ~n426 & n30112;
  assign n30114 = ~n292 & n30113;
  assign n30115 = ~n102 & n30114;
  assign n30116 = ~n422 & n30115;
  assign n30117 = ~n531 & n30116;
  assign n30118 = ~n29946 & n30117;
  assign n30119 = n29946 & ~n30117;
  assign n30120 = ~n30099 & ~n30119;
  assign n30121 = ~n30118 & n30120;
  assign n30122 = ~n30099 & ~n30121;
  assign n30123 = ~n30119 & ~n30121;
  assign n30124 = ~n30118 & n30123;
  assign n30125 = ~n30122 & ~n30124;
  assign n30126 = n75 & ~n23642;
  assign n30127 = n3020 & n22344;
  assign n30128 = n3023 & n22350;
  assign n30129 = n3028 & n22347;
  assign n30130 = ~n30128 & ~n30129;
  assign n30131 = ~n30127 & n30130;
  assign n30132 = ~n30126 & n30131;
  assign n30133 = ~n30125 & ~n30132;
  assign n30134 = ~n30125 & ~n30133;
  assign n30135 = ~n30132 & ~n30133;
  assign n30136 = ~n30134 & ~n30135;
  assign n30137 = n3457 & n22335;
  assign n30138 = n3542 & n22341;
  assign n30139 = n3606 & n22338;
  assign n30140 = ~n30138 & ~n30139;
  assign n30141 = ~n30137 & n30140;
  assign n30142 = ~n3368 & n30141;
  assign n30143 = n24167 & n30141;
  assign n30144 = ~n30142 & ~n30143;
  assign n30145 =  a[29]  & ~n30144;
  assign n30146 = ~ a[29]  & n30144;
  assign n30147 = ~n30145 & ~n30146;
  assign n30148 = ~n30136 & ~n30147;
  assign n30149 = n30136 & n30147;
  assign n30150 = ~n30148 & ~n30149;
  assign n30151 = ~n30098 & n30150;
  assign n30152 = n30098 & ~n30150;
  assign n30153 = ~n30151 & ~n30152;
  assign n30154 = n3884 & n22326;
  assign n30155 = n3967 & n22332;
  assign n30156 = n4046 & n22329;
  assign n30157 = ~n30155 & ~n30156;
  assign n30158 = ~n30154 & n30157;
  assign n30159 = n4050 & ~n24616;
  assign n30160 = n30158 & ~n30159;
  assign n30161 =  a[26]  & ~n30160;
  assign n30162 =  a[26]  & ~n30161;
  assign n30163 = ~n30160 & ~n30161;
  assign n30164 = ~n30162 & ~n30163;
  assign n30165 = n30153 & ~n30164;
  assign n30166 = n30153 & ~n30165;
  assign n30167 = ~n30164 & ~n30165;
  assign n30168 = ~n30166 & ~n30167;
  assign n30169 = ~n29972 & ~n29986;
  assign n30170 = n30168 & n30169;
  assign n30171 = ~n30168 & ~n30169;
  assign n30172 = ~n30170 & ~n30171;
  assign n30173 = n4694 & n22312;
  assign n30174 = n4533 & n22323;
  assign n30175 = n4604 & n22320;
  assign n30176 = ~n30174 & ~n30175;
  assign n30177 = ~n30173 & n30176;
  assign n30178 = n4536 & ~n25315;
  assign n30179 = n30177 & ~n30178;
  assign n30180 =  a[23]  & ~n30179;
  assign n30181 =  a[23]  & ~n30180;
  assign n30182 = ~n30179 & ~n30180;
  assign n30183 = ~n30181 & ~n30182;
  assign n30184 = n30172 & ~n30183;
  assign n30185 = n30172 & ~n30184;
  assign n30186 = ~n30183 & ~n30184;
  assign n30187 = ~n30185 & ~n30186;
  assign n30188 = ~n29992 & ~n30005;
  assign n30189 = n30187 & n30188;
  assign n30190 = ~n30187 & ~n30188;
  assign n30191 = ~n30189 & ~n30190;
  assign n30192 = n5496 & n26063;
  assign n30193 = n4935 & n22315;
  assign n30194 = n5407 & n22309;
  assign n30195 = ~n30193 & ~n30194;
  assign n30196 = ~n30192 & n30195;
  assign n30197 = n4938 & ~n26604;
  assign n30198 = n30196 & ~n30197;
  assign n30199 =  a[20]  & ~n30198;
  assign n30200 =  a[20]  & ~n30199;
  assign n30201 = ~n30198 & ~n30199;
  assign n30202 = ~n30200 & ~n30201;
  assign n30203 = n30191 & ~n30202;
  assign n30204 = n30191 & ~n30203;
  assign n30205 = ~n30202 & ~n30203;
  assign n30206 = ~n30204 & ~n30205;
  assign n30207 = ~n30011 & ~n30024;
  assign n30208 = n30206 & n30207;
  assign n30209 = ~n30206 & ~n30207;
  assign n30210 = ~n30208 & ~n30209;
  assign n30211 = n6233 & n26890;
  assign n30212 = n5663 & n26066;
  assign n30213 = n5939 & n26060;
  assign n30214 = ~n30212 & ~n30213;
  assign n30215 = ~n30211 & n30214;
  assign n30216 = n5666 & ~n26904;
  assign n30217 = n30215 & ~n30216;
  assign n30218 =  a[17]  & ~n30217;
  assign n30219 =  a[17]  & ~n30218;
  assign n30220 = ~n30217 & ~n30218;
  assign n30221 = ~n30219 & ~n30220;
  assign n30222 = n30210 & ~n30221;
  assign n30223 = n30210 & ~n30222;
  assign n30224 = ~n30221 & ~n30222;
  assign n30225 = ~n30223 & ~n30224;
  assign n30226 = ~n30030 & ~n30043;
  assign n30227 = n30225 & n30226;
  assign n30228 = ~n30225 & ~n30226;
  assign n30229 = ~n30227 & ~n30228;
  assign n30230 = n7101 & n27698;
  assign n30231 = n6402 & n27173;
  assign n30232 = n6951 & n27442;
  assign n30233 = ~n30231 & ~n30232;
  assign n30234 = ~n30230 & n30233;
  assign n30235 = n6397 & ~n27713;
  assign n30236 = n30234 & ~n30235;
  assign n30237 =  a[14]  & ~n30236;
  assign n30238 =  a[14]  & ~n30237;
  assign n30239 = ~n30236 & ~n30237;
  assign n30240 = ~n30238 & ~n30239;
  assign n30241 = n30229 & ~n30240;
  assign n30242 = n30229 & ~n30241;
  assign n30243 = ~n30240 & ~n30241;
  assign n30244 = ~n30242 & ~n30243;
  assign n30245 = ~n30048 & ~n30063;
  assign n30246 = ~n14424 & ~n28208;
  assign n30247 = n7291 & n27964;
  assign n30248 = ~n30246 & ~n30247;
  assign n30249 = ~n7294 & n30248;
  assign n30250 = n28221 & n30248;
  assign n30251 = ~n30249 & ~n30250;
  assign n30252 =  a[11]  & ~n30251;
  assign n30253 = ~ a[11]  & n30251;
  assign n30254 = ~n30252 & ~n30253;
  assign n30255 = ~n30245 & ~n30254;
  assign n30256 = n30245 & n30254;
  assign n30257 = ~n30255 & ~n30256;
  assign n30258 = ~n30244 & n30257;
  assign n30259 = ~n30244 & ~n30258;
  assign n30260 = n30257 & ~n30258;
  assign n30261 = ~n30259 & ~n30260;
  assign n30262 = ~n30069 & ~n30082;
  assign n30263 = n30261 & n30262;
  assign n30264 = ~n30261 & ~n30262;
  assign n30265 = ~n30263 & ~n30264;
  assign n30266 = ~n30087 & ~n30093;
  assign n30267 = ~n30265 & n30266;
  assign n30268 = n30265 & ~n30266;
  assign n30269 = ~n30267 & ~n30268;
  assign n30270 = n29921 & n30094;
  assign n30271 = n30269 & n30270;
  assign n30272 = ~n30269 & ~n30270;
  assign  result[15]  = ~n30271 & ~n30272;
  assign n30274 = ~n30264 & ~n30268;
  assign n30275 = ~n30255 & ~n30258;
  assign n30276 = ~n30133 & ~n30148;
  assign n30277 = n75 & n24142;
  assign n30278 = n3020 & n22341;
  assign n30279 = n3023 & n22347;
  assign n30280 = n3028 & n22344;
  assign n30281 = ~n30279 & ~n30280;
  assign n30282 = ~n30278 & n30281;
  assign n30283 = ~n30277 & n30282;
  assign n30284 = ~n14426 & ~n28208;
  assign n30285 =  a[11]  & ~n30284;
  assign n30286 = ~ a[11]  & n30284;
  assign n30287 = ~n30285 & ~n30286;
  assign n30288 = n675 & n2174;
  assign n30289 = n5038 & n30288;
  assign n30290 = n2808 & n30289;
  assign n30291 = n5019 & n30290;
  assign n30292 = n1407 & n30291;
  assign n30293 = n3510 & n30292;
  assign n30294 = n241 & n30293;
  assign n30295 = n1435 & n30294;
  assign n30296 = n1576 & n30295;
  assign n30297 = n1252 & n30296;
  assign n30298 = n3886 & n30297;
  assign n30299 = n590 & n30298;
  assign n30300 = ~n242 & n30299;
  assign n30301 = ~n435 & n30300;
  assign n30302 = ~n532 & n30301;
  assign n30303 = ~n363 & n30302;
  assign n30304 = n29946 & n30303;
  assign n30305 = ~n29946 & ~n30303;
  assign n30306 = ~n30304 & ~n30305;
  assign n30307 = n30287 & n30306;
  assign n30308 = ~n30287 & ~n30306;
  assign n30309 = ~n30307 & ~n30308;
  assign n30310 = ~n30283 & n30309;
  assign n30311 = n30309 & ~n30310;
  assign n30312 = ~n30283 & ~n30310;
  assign n30313 = ~n30311 & ~n30312;
  assign n30314 = ~n30123 & ~n30313;
  assign n30315 = ~n30313 & ~n30314;
  assign n30316 = ~n30123 & ~n30314;
  assign n30317 = ~n30315 & ~n30316;
  assign n30318 = ~n30276 & ~n30317;
  assign n30319 = ~n30276 & ~n30318;
  assign n30320 = ~n30317 & ~n30318;
  assign n30321 = ~n30319 & ~n30320;
  assign n30322 = n3457 & n22332;
  assign n30323 = n3542 & n22338;
  assign n30324 = n3606 & n22335;
  assign n30325 = ~n30323 & ~n30324;
  assign n30326 = ~n30322 & n30325;
  assign n30327 = n3368 & n22542;
  assign n30328 = n30326 & ~n30327;
  assign n30329 =  a[29]  & ~n30328;
  assign n30330 =  a[29]  & ~n30329;
  assign n30331 = ~n30328 & ~n30329;
  assign n30332 = ~n30330 & ~n30331;
  assign n30333 = ~n30321 & ~n30332;
  assign n30334 = ~n30321 & ~n30333;
  assign n30335 = ~n30332 & ~n30333;
  assign n30336 = ~n30334 & ~n30335;
  assign n30337 = n3884 & n22323;
  assign n30338 = n3967 & n22329;
  assign n30339 = n4046 & n22326;
  assign n30340 = ~n30338 & ~n30339;
  assign n30341 = ~n30337 & n30340;
  assign n30342 = n4050 & n24599;
  assign n30343 = n30341 & ~n30342;
  assign n30344 =  a[26]  & ~n30343;
  assign n30345 =  a[26]  & ~n30344;
  assign n30346 = ~n30343 & ~n30344;
  assign n30347 = ~n30345 & ~n30346;
  assign n30348 = ~n30336 & ~n30347;
  assign n30349 = ~n30336 & ~n30348;
  assign n30350 = ~n30347 & ~n30348;
  assign n30351 = ~n30349 & ~n30350;
  assign n30352 = ~n30151 & ~n30165;
  assign n30353 = n30351 & n30352;
  assign n30354 = ~n30351 & ~n30352;
  assign n30355 = ~n30353 & ~n30354;
  assign n30356 = n4694 & n22315;
  assign n30357 = n4533 & n22320;
  assign n30358 = n4604 & n22312;
  assign n30359 = ~n30357 & ~n30358;
  assign n30360 = ~n30356 & n30359;
  assign n30361 = n4536 & n25294;
  assign n30362 = n30360 & ~n30361;
  assign n30363 =  a[23]  & ~n30362;
  assign n30364 =  a[23]  & ~n30363;
  assign n30365 = ~n30362 & ~n30363;
  assign n30366 = ~n30364 & ~n30365;
  assign n30367 = n30355 & ~n30366;
  assign n30368 = n30355 & ~n30367;
  assign n30369 = ~n30366 & ~n30367;
  assign n30370 = ~n30368 & ~n30369;
  assign n30371 = ~n30171 & ~n30184;
  assign n30372 = n30370 & n30371;
  assign n30373 = ~n30370 & ~n30371;
  assign n30374 = ~n30372 & ~n30373;
  assign n30375 = ~n30190 & ~n30203;
  assign n30376 = n5496 & n26066;
  assign n30377 = n4935 & n22309;
  assign n30378 = n5407 & n26063;
  assign n30379 = ~n30377 & ~n30378;
  assign n30380 = ~n30376 & n30379;
  assign n30381 = n4938 & ~n26624;
  assign n30382 = n30380 & ~n30381;
  assign n30383 =  a[20]  & ~n30382;
  assign n30384 =  a[20]  & ~n30383;
  assign n30385 = ~n30382 & ~n30383;
  assign n30386 = ~n30384 & ~n30385;
  assign n30387 = ~n30375 & ~n30386;
  assign n30388 = ~n30375 & ~n30387;
  assign n30389 = ~n30386 & ~n30387;
  assign n30390 = ~n30388 & ~n30389;
  assign n30391 = ~n30374 & n30390;
  assign n30392 = n30374 & ~n30390;
  assign n30393 = ~n30391 & ~n30392;
  assign n30394 = n6233 & n27173;
  assign n30395 = n5663 & n26060;
  assign n30396 = n5939 & n26890;
  assign n30397 = ~n30395 & ~n30396;
  assign n30398 = ~n30394 & n30397;
  assign n30399 = n5666 & n27185;
  assign n30400 = n30398 & ~n30399;
  assign n30401 =  a[17]  & ~n30400;
  assign n30402 =  a[17]  & ~n30401;
  assign n30403 = ~n30400 & ~n30401;
  assign n30404 = ~n30402 & ~n30403;
  assign n30405 = n30393 & ~n30404;
  assign n30406 = n30393 & ~n30405;
  assign n30407 = ~n30404 & ~n30405;
  assign n30408 = ~n30406 & ~n30407;
  assign n30409 = ~n30209 & ~n30222;
  assign n30410 = n30408 & n30409;
  assign n30411 = ~n30408 & ~n30409;
  assign n30412 = ~n30410 & ~n30411;
  assign n30413 = ~n30228 & ~n30241;
  assign n30414 = n7101 & n27964;
  assign n30415 = n6402 & n27442;
  assign n30416 = n6951 & n27698;
  assign n30417 = ~n30415 & ~n30416;
  assign n30418 = ~n30414 & n30417;
  assign n30419 = n6397 & n27976;
  assign n30420 = n30418 & ~n30419;
  assign n30421 =  a[14]  & ~n30420;
  assign n30422 =  a[14]  & ~n30421;
  assign n30423 = ~n30420 & ~n30421;
  assign n30424 = ~n30422 & ~n30423;
  assign n30425 = ~n30413 & ~n30424;
  assign n30426 = ~n30413 & ~n30425;
  assign n30427 = ~n30424 & ~n30425;
  assign n30428 = ~n30426 & ~n30427;
  assign n30429 = ~n30412 & n30428;
  assign n30430 = n30412 & ~n30428;
  assign n30431 = ~n30429 & ~n30430;
  assign n30432 = ~n30275 & n30431;
  assign n30433 = n30275 & ~n30431;
  assign n30434 = ~n30432 & ~n30433;
  assign n30435 = ~n30274 & n30434;
  assign n30436 = n30274 & ~n30434;
  assign n30437 = ~n30435 & ~n30436;
  assign n30438 = ~n30271 & ~n30437;
  assign n30439 = n30271 & n30437;
  assign  result[16]  = ~n30438 & ~n30439;
  assign n30441 = ~n30318 & ~n30333;
  assign n30442 = n75 & ~n24188;
  assign n30443 = n3020 & n22338;
  assign n30444 = n3023 & n22344;
  assign n30445 = n3028 & n22341;
  assign n30446 = ~n30444 & ~n30445;
  assign n30447 = ~n30443 & n30446;
  assign n30448 = ~n30442 & n30447;
  assign n30449 = ~n30305 & ~n30307;
  assign n30450 = n1499 & n2059;
  assign n30451 = n778 & n30450;
  assign n30452 = n3128 & n30451;
  assign n30453 = n12977 & n30452;
  assign n30454 = n27789 & n30453;
  assign n30455 = n13458 & n30454;
  assign n30456 = n15324 & n30455;
  assign n30457 = n28294 & n30456;
  assign n30458 = n1380 & n30457;
  assign n30459 = n810 & n30458;
  assign n30460 = ~n469 & n30459;
  assign n30461 = ~n746 & n30460;
  assign n30462 = ~n1102 & n30461;
  assign n30463 = ~n396 & n30462;
  assign n30464 = ~n470 & n30463;
  assign n30465 = ~n30449 & n30464;
  assign n30466 = n30449 & ~n30464;
  assign n30467 = ~n30465 & ~n30466;
  assign n30468 = ~n30448 & n30467;
  assign n30469 = ~n30448 & ~n30468;
  assign n30470 = n30467 & ~n30468;
  assign n30471 = ~n30469 & ~n30470;
  assign n30472 = ~n30310 & ~n30314;
  assign n30473 = n30471 & n30472;
  assign n30474 = ~n30471 & ~n30472;
  assign n30475 = ~n30473 & ~n30474;
  assign n30476 = n3457 & n22329;
  assign n30477 = n3542 & n22335;
  assign n30478 = n3606 & n22332;
  assign n30479 = ~n30477 & ~n30478;
  assign n30480 = ~n30476 & n30479;
  assign n30481 = ~n3368 & n30480;
  assign n30482 = n24633 & n30480;
  assign n30483 = ~n30481 & ~n30482;
  assign n30484 =  a[29]  & ~n30483;
  assign n30485 = ~ a[29]  & n30483;
  assign n30486 = ~n30484 & ~n30485;
  assign n30487 = n30475 & ~n30486;
  assign n30488 = ~n30475 & n30486;
  assign n30489 = ~n30487 & ~n30488;
  assign n30490 = ~n30441 & n30489;
  assign n30491 = n30441 & ~n30489;
  assign n30492 = ~n30490 & ~n30491;
  assign n30493 = n3884 & n22320;
  assign n30494 = n3967 & n22326;
  assign n30495 = n4046 & n22323;
  assign n30496 = ~n30494 & ~n30495;
  assign n30497 = ~n30493 & n30496;
  assign n30498 = n4050 & ~n25270;
  assign n30499 = n30497 & ~n30498;
  assign n30500 =  a[26]  & ~n30499;
  assign n30501 =  a[26]  & ~n30500;
  assign n30502 = ~n30499 & ~n30500;
  assign n30503 = ~n30501 & ~n30502;
  assign n30504 = n30492 & ~n30503;
  assign n30505 = n30492 & ~n30504;
  assign n30506 = ~n30503 & ~n30504;
  assign n30507 = ~n30505 & ~n30506;
  assign n30508 = ~n30348 & ~n30354;
  assign n30509 = n30507 & n30508;
  assign n30510 = ~n30507 & ~n30508;
  assign n30511 = ~n30509 & ~n30510;
  assign n30512 = n4694 & n22309;
  assign n30513 = n4533 & n22312;
  assign n30514 = n4604 & n22315;
  assign n30515 = ~n30513 & ~n30514;
  assign n30516 = ~n30512 & n30515;
  assign n30517 = n4536 & ~n22529;
  assign n30518 = n30516 & ~n30517;
  assign n30519 =  a[23]  & ~n30518;
  assign n30520 =  a[23]  & ~n30519;
  assign n30521 = ~n30518 & ~n30519;
  assign n30522 = ~n30520 & ~n30521;
  assign n30523 = n30511 & ~n30522;
  assign n30524 = n30511 & ~n30523;
  assign n30525 = ~n30522 & ~n30523;
  assign n30526 = ~n30524 & ~n30525;
  assign n30527 = ~n30367 & ~n30373;
  assign n30528 = n30526 & n30527;
  assign n30529 = ~n30526 & ~n30527;
  assign n30530 = ~n30528 & ~n30529;
  assign n30531 = n5496 & n26060;
  assign n30532 = n4935 & n26063;
  assign n30533 = n5407 & n26066;
  assign n30534 = ~n30532 & ~n30533;
  assign n30535 = ~n30531 & n30534;
  assign n30536 = n4938 & ~n26088;
  assign n30537 = n30535 & ~n30536;
  assign n30538 =  a[20]  & ~n30537;
  assign n30539 =  a[20]  & ~n30538;
  assign n30540 = ~n30537 & ~n30538;
  assign n30541 = ~n30539 & ~n30540;
  assign n30542 = n30530 & ~n30541;
  assign n30543 = n30530 & ~n30542;
  assign n30544 = ~n30541 & ~n30542;
  assign n30545 = ~n30543 & ~n30544;
  assign n30546 = ~n30387 & ~n30392;
  assign n30547 = ~n30545 & ~n30546;
  assign n30548 = ~n30545 & ~n30547;
  assign n30549 = ~n30546 & ~n30547;
  assign n30550 = ~n30548 & ~n30549;
  assign n30551 = n6233 & n27442;
  assign n30552 = n5663 & n26890;
  assign n30553 = n5939 & n27173;
  assign n30554 = ~n30552 & ~n30553;
  assign n30555 = ~n30551 & n30554;
  assign n30556 = n5666 & n27455;
  assign n30557 = n30555 & ~n30556;
  assign n30558 =  a[17]  & ~n30557;
  assign n30559 =  a[17]  & ~n30558;
  assign n30560 = ~n30557 & ~n30558;
  assign n30561 = ~n30559 & ~n30560;
  assign n30562 = ~n30550 & ~n30561;
  assign n30563 = ~n30550 & ~n30562;
  assign n30564 = ~n30561 & ~n30562;
  assign n30565 = ~n30563 & ~n30564;
  assign n30566 = ~n30405 & ~n30411;
  assign n30567 = n30565 & n30566;
  assign n30568 = ~n30565 & ~n30566;
  assign n30569 = ~n30567 & ~n30568;
  assign n30570 = n7101 & ~n28208;
  assign n30571 = n6402 & n27698;
  assign n30572 = n6951 & n27964;
  assign n30573 = ~n30571 & ~n30572;
  assign n30574 = ~n30570 & n30573;
  assign n30575 = n6397 & ~n28223;
  assign n30576 = n30574 & ~n30575;
  assign n30577 =  a[14]  & ~n30576;
  assign n30578 =  a[14]  & ~n30577;
  assign n30579 = ~n30576 & ~n30577;
  assign n30580 = ~n30578 & ~n30579;
  assign n30581 = n30569 & ~n30580;
  assign n30582 = n30569 & ~n30581;
  assign n30583 = ~n30580 & ~n30581;
  assign n30584 = ~n30582 & ~n30583;
  assign n30585 = ~n30425 & ~n30430;
  assign n30586 = ~n30584 & ~n30585;
  assign n30587 = ~n30584 & ~n30586;
  assign n30588 = ~n30585 & ~n30586;
  assign n30589 = ~n30587 & ~n30588;
  assign n30590 = ~n30432 & ~n30435;
  assign n30591 = n30589 & n30590;
  assign n30592 = ~n30589 & ~n30590;
  assign n30593 = ~n30591 & ~n30592;
  assign n30594 = ~n30439 & n30593;
  assign n30595 = n30439 & ~n30593;
  assign  result[17]  = n30594 | n30595;
  assign n30597 = n30439 & n30593;
  assign n30598 = n75 & ~n24167;
  assign n30599 = n3020 & n22335;
  assign n30600 = n3023 & n22341;
  assign n30601 = n3028 & n22338;
  assign n30602 = ~n30600 & ~n30601;
  assign n30603 = ~n30599 & n30602;
  assign n30604 = ~n30598 & n30603;
  assign n30605 = n694 & n2176;
  assign n30606 = n6084 & n30605;
  assign n30607 = n3108 & n30606;
  assign n30608 = n12710 & n30607;
  assign n30609 = n13123 & n30608;
  assign n30610 = n3386 & n30609;
  assign n30611 = n2500 & n30610;
  assign n30612 = n5209 & n30611;
  assign n30613 = n2739 & n30612;
  assign n30614 = ~n558 & n30613;
  assign n30615 = ~n1102 & n30614;
  assign n30616 = ~n155 & n30615;
  assign n30617 = ~n248 & n30616;
  assign n30618 = ~n357 & n30617;
  assign n30619 = ~n205 & n30618;
  assign n30620 = ~n436 & n30619;
  assign n30621 = ~n81 & n30620;
  assign n30622 = ~n30464 & n30621;
  assign n30623 = n30464 & ~n30621;
  assign n30624 = ~n30604 & ~n30623;
  assign n30625 = ~n30622 & n30624;
  assign n30626 = ~n30604 & ~n30625;
  assign n30627 = ~n30623 & ~n30625;
  assign n30628 = ~n30622 & n30627;
  assign n30629 = ~n30626 & ~n30628;
  assign n30630 = ~n30465 & ~n30468;
  assign n30631 = n30629 & n30630;
  assign n30632 = ~n30629 & ~n30630;
  assign n30633 = ~n30631 & ~n30632;
  assign n30634 = ~n30474 & ~n30487;
  assign n30635 = ~n30633 & n30634;
  assign n30636 = n30633 & ~n30634;
  assign n30637 = ~n30635 & ~n30636;
  assign n30638 = n3457 & n22326;
  assign n30639 = n3542 & n22332;
  assign n30640 = n3606 & n22329;
  assign n30641 = ~n30639 & ~n30640;
  assign n30642 = ~n30638 & n30641;
  assign n30643 = n3368 & ~n24616;
  assign n30644 = n30642 & ~n30643;
  assign n30645 =  a[29]  & ~n30644;
  assign n30646 =  a[29]  & ~n30645;
  assign n30647 = ~n30644 & ~n30645;
  assign n30648 = ~n30646 & ~n30647;
  assign n30649 = n30637 & ~n30648;
  assign n30650 = n30637 & ~n30649;
  assign n30651 = ~n30648 & ~n30649;
  assign n30652 = ~n30650 & ~n30651;
  assign n30653 = n3884 & n22312;
  assign n30654 = n3967 & n22323;
  assign n30655 = n4046 & n22320;
  assign n30656 = ~n30654 & ~n30655;
  assign n30657 = ~n30653 & n30656;
  assign n30658 = n4050 & ~n25315;
  assign n30659 = n30657 & ~n30658;
  assign n30660 =  a[26]  & ~n30659;
  assign n30661 =  a[26]  & ~n30660;
  assign n30662 = ~n30659 & ~n30660;
  assign n30663 = ~n30661 & ~n30662;
  assign n30664 = ~n30652 & ~n30663;
  assign n30665 = ~n30652 & ~n30664;
  assign n30666 = ~n30663 & ~n30664;
  assign n30667 = ~n30665 & ~n30666;
  assign n30668 = ~n30490 & ~n30504;
  assign n30669 = n30667 & n30668;
  assign n30670 = ~n30667 & ~n30668;
  assign n30671 = ~n30669 & ~n30670;
  assign n30672 = n4694 & n26063;
  assign n30673 = n4533 & n22315;
  assign n30674 = n4604 & n22309;
  assign n30675 = ~n30673 & ~n30674;
  assign n30676 = ~n30672 & n30675;
  assign n30677 = n4536 & ~n26604;
  assign n30678 = n30676 & ~n30677;
  assign n30679 =  a[23]  & ~n30678;
  assign n30680 =  a[23]  & ~n30679;
  assign n30681 = ~n30678 & ~n30679;
  assign n30682 = ~n30680 & ~n30681;
  assign n30683 = n30671 & ~n30682;
  assign n30684 = n30671 & ~n30683;
  assign n30685 = ~n30682 & ~n30683;
  assign n30686 = ~n30684 & ~n30685;
  assign n30687 = ~n30510 & ~n30523;
  assign n30688 = n30686 & n30687;
  assign n30689 = ~n30686 & ~n30687;
  assign n30690 = ~n30688 & ~n30689;
  assign n30691 = n5496 & n26890;
  assign n30692 = n4935 & n26066;
  assign n30693 = n5407 & n26060;
  assign n30694 = ~n30692 & ~n30693;
  assign n30695 = ~n30691 & n30694;
  assign n30696 = n4938 & ~n26904;
  assign n30697 = n30695 & ~n30696;
  assign n30698 =  a[20]  & ~n30697;
  assign n30699 =  a[20]  & ~n30698;
  assign n30700 = ~n30697 & ~n30698;
  assign n30701 = ~n30699 & ~n30700;
  assign n30702 = n30690 & ~n30701;
  assign n30703 = n30690 & ~n30702;
  assign n30704 = ~n30701 & ~n30702;
  assign n30705 = ~n30703 & ~n30704;
  assign n30706 = ~n30529 & ~n30542;
  assign n30707 = n30705 & n30706;
  assign n30708 = ~n30705 & ~n30706;
  assign n30709 = ~n30707 & ~n30708;
  assign n30710 = n6233 & n27698;
  assign n30711 = n5663 & n27173;
  assign n30712 = n5939 & n27442;
  assign n30713 = ~n30711 & ~n30712;
  assign n30714 = ~n30710 & n30713;
  assign n30715 = n5666 & ~n27713;
  assign n30716 = n30714 & ~n30715;
  assign n30717 =  a[17]  & ~n30716;
  assign n30718 =  a[17]  & ~n30717;
  assign n30719 = ~n30716 & ~n30717;
  assign n30720 = ~n30718 & ~n30719;
  assign n30721 = n30709 & ~n30720;
  assign n30722 = n30709 & ~n30721;
  assign n30723 = ~n30720 & ~n30721;
  assign n30724 = ~n30722 & ~n30723;
  assign n30725 = ~n30547 & ~n30562;
  assign n30726 = ~n13845 & ~n28208;
  assign n30727 = n6402 & n27964;
  assign n30728 = ~n30726 & ~n30727;
  assign n30729 = ~n6397 & n30728;
  assign n30730 = n28221 & n30728;
  assign n30731 = ~n30729 & ~n30730;
  assign n30732 =  a[14]  & ~n30731;
  assign n30733 = ~ a[14]  & n30731;
  assign n30734 = ~n30732 & ~n30733;
  assign n30735 = ~n30725 & ~n30734;
  assign n30736 = n30725 & n30734;
  assign n30737 = ~n30735 & ~n30736;
  assign n30738 = ~n30724 & n30737;
  assign n30739 = ~n30724 & ~n30738;
  assign n30740 = n30737 & ~n30738;
  assign n30741 = ~n30739 & ~n30740;
  assign n30742 = ~n30568 & ~n30581;
  assign n30743 = n30741 & n30742;
  assign n30744 = ~n30741 & ~n30742;
  assign n30745 = ~n30743 & ~n30744;
  assign n30746 = ~n30586 & ~n30592;
  assign n30747 = ~n30745 & n30746;
  assign n30748 = n30745 & ~n30746;
  assign n30749 = ~n30747 & ~n30748;
  assign n30750 = n30597 & n30749;
  assign n30751 = ~n30597 & ~n30749;
  assign  result[18]  = ~n30750 & ~n30751;
  assign n30753 = ~n30744 & ~n30748;
  assign n30754 = ~n30735 & ~n30738;
  assign n30755 = n75 & n22542;
  assign n30756 = n3020 & n22332;
  assign n30757 = n3023 & n22338;
  assign n30758 = n3028 & n22335;
  assign n30759 = ~n30757 & ~n30758;
  assign n30760 = ~n30756 & n30759;
  assign n30761 = ~n30755 & n30760;
  assign n30762 = ~n13847 & ~n28208;
  assign n30763 =  a[14]  & ~n30762;
  assign n30764 = ~ a[14]  & n30762;
  assign n30765 = ~n30763 & ~n30764;
  assign n30766 = n2537 & n3045;
  assign n30767 = n14482 & n30766;
  assign n30768 = n1894 & n30767;
  assign n30769 = n14202 & n30768;
  assign n30770 = n6714 & n30769;
  assign n30771 = n1291 & n30770;
  assign n30772 = n976 & n30771;
  assign n30773 = n1139 & n30772;
  assign n30774 = n2219 & n30773;
  assign n30775 = ~n357 & n30774;
  assign n30776 = ~n326 & n30775;
  assign n30777 = ~n452 & n30776;
  assign n30778 = n30464 & n30777;
  assign n30779 = ~n30464 & ~n30777;
  assign n30780 = ~n30778 & ~n30779;
  assign n30781 = n30765 & n30780;
  assign n30782 = ~n30765 & ~n30780;
  assign n30783 = ~n30781 & ~n30782;
  assign n30784 = ~n30627 & n30783;
  assign n30785 = n30627 & ~n30783;
  assign n30786 = ~n30784 & ~n30785;
  assign n30787 = ~n30761 & n30786;
  assign n30788 = n30786 & ~n30787;
  assign n30789 = ~n30761 & ~n30787;
  assign n30790 = ~n30788 & ~n30789;
  assign n30791 = n3457 & n22323;
  assign n30792 = n3542 & n22329;
  assign n30793 = n3606 & n22326;
  assign n30794 = ~n30792 & ~n30793;
  assign n30795 = ~n30791 & n30794;
  assign n30796 = n3368 & n24599;
  assign n30797 = n30795 & ~n30796;
  assign n30798 =  a[29]  & ~n30797;
  assign n30799 =  a[29]  & ~n30798;
  assign n30800 = ~n30797 & ~n30798;
  assign n30801 = ~n30799 & ~n30800;
  assign n30802 = ~n30790 & ~n30801;
  assign n30803 = ~n30790 & ~n30802;
  assign n30804 = ~n30801 & ~n30802;
  assign n30805 = ~n30803 & ~n30804;
  assign n30806 = ~n30632 & ~n30636;
  assign n30807 = n30805 & n30806;
  assign n30808 = ~n30805 & ~n30806;
  assign n30809 = ~n30807 & ~n30808;
  assign n30810 = n3884 & n22315;
  assign n30811 = n3967 & n22320;
  assign n30812 = n4046 & n22312;
  assign n30813 = ~n30811 & ~n30812;
  assign n30814 = ~n30810 & n30813;
  assign n30815 = n4050 & n25294;
  assign n30816 = n30814 & ~n30815;
  assign n30817 =  a[26]  & ~n30816;
  assign n30818 =  a[26]  & ~n30817;
  assign n30819 = ~n30816 & ~n30817;
  assign n30820 = ~n30818 & ~n30819;
  assign n30821 = n30809 & ~n30820;
  assign n30822 = n30809 & ~n30821;
  assign n30823 = ~n30820 & ~n30821;
  assign n30824 = ~n30822 & ~n30823;
  assign n30825 = ~n30649 & ~n30664;
  assign n30826 = n30824 & n30825;
  assign n30827 = ~n30824 & ~n30825;
  assign n30828 = ~n30826 & ~n30827;
  assign n30829 = ~n30670 & ~n30683;
  assign n30830 = n4694 & n26066;
  assign n30831 = n4533 & n22309;
  assign n30832 = n4604 & n26063;
  assign n30833 = ~n30831 & ~n30832;
  assign n30834 = ~n30830 & n30833;
  assign n30835 = n4536 & ~n26624;
  assign n30836 = n30834 & ~n30835;
  assign n30837 =  a[23]  & ~n30836;
  assign n30838 =  a[23]  & ~n30837;
  assign n30839 = ~n30836 & ~n30837;
  assign n30840 = ~n30838 & ~n30839;
  assign n30841 = ~n30829 & ~n30840;
  assign n30842 = ~n30829 & ~n30841;
  assign n30843 = ~n30840 & ~n30841;
  assign n30844 = ~n30842 & ~n30843;
  assign n30845 = ~n30828 & n30844;
  assign n30846 = n30828 & ~n30844;
  assign n30847 = ~n30845 & ~n30846;
  assign n30848 = n5496 & n27173;
  assign n30849 = n4935 & n26060;
  assign n30850 = n5407 & n26890;
  assign n30851 = ~n30849 & ~n30850;
  assign n30852 = ~n30848 & n30851;
  assign n30853 = n4938 & n27185;
  assign n30854 = n30852 & ~n30853;
  assign n30855 =  a[20]  & ~n30854;
  assign n30856 =  a[20]  & ~n30855;
  assign n30857 = ~n30854 & ~n30855;
  assign n30858 = ~n30856 & ~n30857;
  assign n30859 = n30847 & ~n30858;
  assign n30860 = n30847 & ~n30859;
  assign n30861 = ~n30858 & ~n30859;
  assign n30862 = ~n30860 & ~n30861;
  assign n30863 = ~n30689 & ~n30702;
  assign n30864 = n30862 & n30863;
  assign n30865 = ~n30862 & ~n30863;
  assign n30866 = ~n30864 & ~n30865;
  assign n30867 = ~n30708 & ~n30721;
  assign n30868 = n6233 & n27964;
  assign n30869 = n5663 & n27442;
  assign n30870 = n5939 & n27698;
  assign n30871 = ~n30869 & ~n30870;
  assign n30872 = ~n30868 & n30871;
  assign n30873 = n5666 & n27976;
  assign n30874 = n30872 & ~n30873;
  assign n30875 =  a[17]  & ~n30874;
  assign n30876 =  a[17]  & ~n30875;
  assign n30877 = ~n30874 & ~n30875;
  assign n30878 = ~n30876 & ~n30877;
  assign n30879 = ~n30867 & ~n30878;
  assign n30880 = ~n30867 & ~n30879;
  assign n30881 = ~n30878 & ~n30879;
  assign n30882 = ~n30880 & ~n30881;
  assign n30883 = ~n30866 & n30882;
  assign n30884 = n30866 & ~n30882;
  assign n30885 = ~n30883 & ~n30884;
  assign n30886 = ~n30754 & n30885;
  assign n30887 = n30754 & ~n30885;
  assign n30888 = ~n30886 & ~n30887;
  assign n30889 = ~n30753 & n30888;
  assign n30890 = n30753 & ~n30888;
  assign n30891 = ~n30889 & ~n30890;
  assign n30892 = ~n30750 & ~n30891;
  assign n30893 = n30750 & n30891;
  assign  result[19]  = ~n30892 & ~n30893;
  assign n30895 = ~n30802 & ~n30808;
  assign n30896 = n75 & ~n24633;
  assign n30897 = n3020 & n22329;
  assign n30898 = n3023 & n22335;
  assign n30899 = n3028 & n22332;
  assign n30900 = ~n30898 & ~n30899;
  assign n30901 = ~n30897 & n30900;
  assign n30902 = ~n30896 & n30901;
  assign n30903 = ~n30779 & ~n30781;
  assign n30904 = n1369 & n3393;
  assign n30905 = n2361 & n30904;
  assign n30906 = n14525 & n30905;
  assign n30907 = n5034 & n30906;
  assign n30908 = n5773 & n30907;
  assign n30909 = n977 & n30908;
  assign n30910 = n491 & n30909;
  assign n30911 = n1183 & n30910;
  assign n30912 = n2346 & n30911;
  assign n30913 = n2697 & n30912;
  assign n30914 = n471 & n30913;
  assign n30915 = n1782 & n30914;
  assign n30916 = ~n224 & n30915;
  assign n30917 = ~n146 & n30916;
  assign n30918 = ~n161 & n30917;
  assign n30919 = ~n358 & n30918;
  assign n30920 = ~n30903 & n30919;
  assign n30921 = n30903 & ~n30919;
  assign n30922 = ~n30920 & ~n30921;
  assign n30923 = ~n30902 & n30922;
  assign n30924 = ~n30902 & ~n30923;
  assign n30925 = n30922 & ~n30923;
  assign n30926 = ~n30924 & ~n30925;
  assign n30927 = ~n30784 & ~n30787;
  assign n30928 = n30926 & n30927;
  assign n30929 = ~n30926 & ~n30927;
  assign n30930 = ~n30928 & ~n30929;
  assign n30931 = n3457 & n22320;
  assign n30932 = n3542 & n22326;
  assign n30933 = n3606 & n22323;
  assign n30934 = ~n30932 & ~n30933;
  assign n30935 = ~n30931 & n30934;
  assign n30936 = ~n3368 & n30935;
  assign n30937 = n25270 & n30935;
  assign n30938 = ~n30936 & ~n30937;
  assign n30939 =  a[29]  & ~n30938;
  assign n30940 = ~ a[29]  & n30938;
  assign n30941 = ~n30939 & ~n30940;
  assign n30942 = n30930 & ~n30941;
  assign n30943 = ~n30930 & n30941;
  assign n30944 = ~n30942 & ~n30943;
  assign n30945 = ~n30895 & n30944;
  assign n30946 = n30895 & ~n30944;
  assign n30947 = ~n30945 & ~n30946;
  assign n30948 = n3884 & n22309;
  assign n30949 = n3967 & n22312;
  assign n30950 = n4046 & n22315;
  assign n30951 = ~n30949 & ~n30950;
  assign n30952 = ~n30948 & n30951;
  assign n30953 = n4050 & ~n22529;
  assign n30954 = n30952 & ~n30953;
  assign n30955 =  a[26]  & ~n30954;
  assign n30956 =  a[26]  & ~n30955;
  assign n30957 = ~n30954 & ~n30955;
  assign n30958 = ~n30956 & ~n30957;
  assign n30959 = n30947 & ~n30958;
  assign n30960 = n30947 & ~n30959;
  assign n30961 = ~n30958 & ~n30959;
  assign n30962 = ~n30960 & ~n30961;
  assign n30963 = ~n30821 & ~n30827;
  assign n30964 = n30962 & n30963;
  assign n30965 = ~n30962 & ~n30963;
  assign n30966 = ~n30964 & ~n30965;
  assign n30967 = n4694 & n26060;
  assign n30968 = n4533 & n26063;
  assign n30969 = n4604 & n26066;
  assign n30970 = ~n30968 & ~n30969;
  assign n30971 = ~n30967 & n30970;
  assign n30972 = n4536 & ~n26088;
  assign n30973 = n30971 & ~n30972;
  assign n30974 =  a[23]  & ~n30973;
  assign n30975 =  a[23]  & ~n30974;
  assign n30976 = ~n30973 & ~n30974;
  assign n30977 = ~n30975 & ~n30976;
  assign n30978 = n30966 & ~n30977;
  assign n30979 = n30966 & ~n30978;
  assign n30980 = ~n30977 & ~n30978;
  assign n30981 = ~n30979 & ~n30980;
  assign n30982 = ~n30841 & ~n30846;
  assign n30983 = ~n30981 & ~n30982;
  assign n30984 = ~n30981 & ~n30983;
  assign n30985 = ~n30982 & ~n30983;
  assign n30986 = ~n30984 & ~n30985;
  assign n30987 = n5496 & n27442;
  assign n30988 = n4935 & n26890;
  assign n30989 = n5407 & n27173;
  assign n30990 = ~n30988 & ~n30989;
  assign n30991 = ~n30987 & n30990;
  assign n30992 = n4938 & n27455;
  assign n30993 = n30991 & ~n30992;
  assign n30994 =  a[20]  & ~n30993;
  assign n30995 =  a[20]  & ~n30994;
  assign n30996 = ~n30993 & ~n30994;
  assign n30997 = ~n30995 & ~n30996;
  assign n30998 = ~n30986 & ~n30997;
  assign n30999 = ~n30986 & ~n30998;
  assign n31000 = ~n30997 & ~n30998;
  assign n31001 = ~n30999 & ~n31000;
  assign n31002 = ~n30859 & ~n30865;
  assign n31003 = n31001 & n31002;
  assign n31004 = ~n31001 & ~n31002;
  assign n31005 = ~n31003 & ~n31004;
  assign n31006 = n6233 & ~n28208;
  assign n31007 = n5663 & n27698;
  assign n31008 = n5939 & n27964;
  assign n31009 = ~n31007 & ~n31008;
  assign n31010 = ~n31006 & n31009;
  assign n31011 = n5666 & ~n28223;
  assign n31012 = n31010 & ~n31011;
  assign n31013 =  a[17]  & ~n31012;
  assign n31014 =  a[17]  & ~n31013;
  assign n31015 = ~n31012 & ~n31013;
  assign n31016 = ~n31014 & ~n31015;
  assign n31017 = n31005 & ~n31016;
  assign n31018 = n31005 & ~n31017;
  assign n31019 = ~n31016 & ~n31017;
  assign n31020 = ~n31018 & ~n31019;
  assign n31021 = ~n30879 & ~n30884;
  assign n31022 = ~n31020 & ~n31021;
  assign n31023 = ~n31020 & ~n31022;
  assign n31024 = ~n31021 & ~n31022;
  assign n31025 = ~n31023 & ~n31024;
  assign n31026 = ~n30886 & ~n30889;
  assign n31027 = n31025 & n31026;
  assign n31028 = ~n31025 & ~n31026;
  assign n31029 = ~n31027 & ~n31028;
  assign n31030 = n30893 & ~n31029;
  assign n31031 = ~n30893 & n31029;
  assign  result[20]  = n31030 | n31031;
  assign n31033 = ~n30929 & ~n30942;
  assign n31034 = ~n30920 & ~n30923;
  assign n31035 = ~n242 & n1253;
  assign n31036 = ~n135 & n31035;
  assign n31037 = n376 & n2026;
  assign n31038 = n31036 & n31037;
  assign n31039 = n2263 & n31038;
  assign n31040 = n5188 & n31039;
  assign n31041 = n13247 & n31040;
  assign n31042 = n1100 & n31041;
  assign n31043 = n2506 & n31042;
  assign n31044 = n1781 & n31043;
  assign n31045 = n3739 & n31044;
  assign n31046 = n1380 & n31045;
  assign n31047 = ~n1306 & n31046;
  assign n31048 = ~n292 & n31047;
  assign n31049 = ~n240 & n31048;
  assign n31050 = ~n225 & n31049;
  assign n31051 = ~n525 & n31050;
  assign n31052 = ~n489 & n31051;
  assign n31053 = n30919 & ~n31052;
  assign n31054 = ~n30919 & n31052;
  assign n31055 = ~n31034 & ~n31054;
  assign n31056 = ~n31053 & n31055;
  assign n31057 = ~n31034 & ~n31056;
  assign n31058 = ~n31054 & ~n31056;
  assign n31059 = ~n31053 & n31058;
  assign n31060 = ~n31057 & ~n31059;
  assign n31061 = n75 & ~n24616;
  assign n31062 = n3020 & n22326;
  assign n31063 = n3023 & n22332;
  assign n31064 = n3028 & n22329;
  assign n31065 = ~n31063 & ~n31064;
  assign n31066 = ~n31062 & n31065;
  assign n31067 = ~n31061 & n31066;
  assign n31068 = ~n31060 & ~n31067;
  assign n31069 = ~n31060 & ~n31068;
  assign n31070 = ~n31067 & ~n31068;
  assign n31071 = ~n31069 & ~n31070;
  assign n31072 = n3457 & n22312;
  assign n31073 = n3542 & n22323;
  assign n31074 = n3606 & n22320;
  assign n31075 = ~n31073 & ~n31074;
  assign n31076 = ~n31072 & n31075;
  assign n31077 = ~n3368 & n31076;
  assign n31078 = n25315 & n31076;
  assign n31079 = ~n31077 & ~n31078;
  assign n31080 =  a[29]  & ~n31079;
  assign n31081 = ~ a[29]  & n31079;
  assign n31082 = ~n31080 & ~n31081;
  assign n31083 = ~n31071 & ~n31082;
  assign n31084 = n31071 & n31082;
  assign n31085 = ~n31083 & ~n31084;
  assign n31086 = ~n31033 & n31085;
  assign n31087 = n31033 & ~n31085;
  assign n31088 = ~n31086 & ~n31087;
  assign n31089 = n3884 & n26063;
  assign n31090 = n3967 & n22315;
  assign n31091 = n4046 & n22309;
  assign n31092 = ~n31090 & ~n31091;
  assign n31093 = ~n31089 & n31092;
  assign n31094 = n4050 & ~n26604;
  assign n31095 = n31093 & ~n31094;
  assign n31096 =  a[26]  & ~n31095;
  assign n31097 =  a[26]  & ~n31096;
  assign n31098 = ~n31095 & ~n31096;
  assign n31099 = ~n31097 & ~n31098;
  assign n31100 = n31088 & ~n31099;
  assign n31101 = n31088 & ~n31100;
  assign n31102 = ~n31099 & ~n31100;
  assign n31103 = ~n31101 & ~n31102;
  assign n31104 = ~n30945 & ~n30959;
  assign n31105 = n31103 & n31104;
  assign n31106 = ~n31103 & ~n31104;
  assign n31107 = ~n31105 & ~n31106;
  assign n31108 = n4694 & n26890;
  assign n31109 = n4533 & n26066;
  assign n31110 = n4604 & n26060;
  assign n31111 = ~n31109 & ~n31110;
  assign n31112 = ~n31108 & n31111;
  assign n31113 = n4536 & ~n26904;
  assign n31114 = n31112 & ~n31113;
  assign n31115 =  a[23]  & ~n31114;
  assign n31116 =  a[23]  & ~n31115;
  assign n31117 = ~n31114 & ~n31115;
  assign n31118 = ~n31116 & ~n31117;
  assign n31119 = n31107 & ~n31118;
  assign n31120 = n31107 & ~n31119;
  assign n31121 = ~n31118 & ~n31119;
  assign n31122 = ~n31120 & ~n31121;
  assign n31123 = ~n30965 & ~n30978;
  assign n31124 = n31122 & n31123;
  assign n31125 = ~n31122 & ~n31123;
  assign n31126 = ~n31124 & ~n31125;
  assign n31127 = n5496 & n27698;
  assign n31128 = n4935 & n27173;
  assign n31129 = n5407 & n27442;
  assign n31130 = ~n31128 & ~n31129;
  assign n31131 = ~n31127 & n31130;
  assign n31132 = n4938 & ~n27713;
  assign n31133 = n31131 & ~n31132;
  assign n31134 =  a[20]  & ~n31133;
  assign n31135 =  a[20]  & ~n31134;
  assign n31136 = ~n31133 & ~n31134;
  assign n31137 = ~n31135 & ~n31136;
  assign n31138 = n31126 & ~n31137;
  assign n31139 = n31126 & ~n31138;
  assign n31140 = ~n31137 & ~n31138;
  assign n31141 = ~n31139 & ~n31140;
  assign n31142 = ~n30983 & ~n30998;
  assign n31143 = ~n13717 & ~n28208;
  assign n31144 = n5663 & n27964;
  assign n31145 = ~n31143 & ~n31144;
  assign n31146 = ~n5666 & n31145;
  assign n31147 = n28221 & n31145;
  assign n31148 = ~n31146 & ~n31147;
  assign n31149 =  a[17]  & ~n31148;
  assign n31150 = ~ a[17]  & n31148;
  assign n31151 = ~n31149 & ~n31150;
  assign n31152 = ~n31142 & ~n31151;
  assign n31153 = n31142 & n31151;
  assign n31154 = ~n31152 & ~n31153;
  assign n31155 = ~n31141 & n31154;
  assign n31156 = ~n31141 & ~n31155;
  assign n31157 = n31154 & ~n31155;
  assign n31158 = ~n31156 & ~n31157;
  assign n31159 = ~n31004 & ~n31017;
  assign n31160 = n31158 & n31159;
  assign n31161 = ~n31158 & ~n31159;
  assign n31162 = ~n31160 & ~n31161;
  assign n31163 = ~n31022 & ~n31028;
  assign n31164 = ~n31162 & n31163;
  assign n31165 = n31162 & ~n31163;
  assign n31166 = ~n31164 & ~n31165;
  assign n31167 = n30893 & n31029;
  assign n31168 = n31166 & n31167;
  assign n31169 = ~n31166 & ~n31167;
  assign  result[21]  = ~n31168 & ~n31169;
  assign n31171 = ~n31161 & ~n31165;
  assign n31172 = ~n31152 & ~n31155;
  assign n31173 = ~n31106 & ~n31119;
  assign n31174 = ~n31086 & ~n31100;
  assign n31175 = n3884 & n26066;
  assign n31176 = n3967 & n22309;
  assign n31177 = n4046 & n26063;
  assign n31178 = ~n31176 & ~n31177;
  assign n31179 = ~n31175 & n31178;
  assign n31180 = n4050 & ~n26624;
  assign n31181 = n31179 & ~n31180;
  assign n31182 =  a[26]  & ~n31181;
  assign n31183 =  a[26]  & ~n31182;
  assign n31184 = ~n31181 & ~n31182;
  assign n31185 = ~n31183 & ~n31184;
  assign n31186 = ~n31174 & ~n31185;
  assign n31187 = ~n31174 & ~n31186;
  assign n31188 = ~n31185 & ~n31186;
  assign n31189 = ~n31187 & ~n31188;
  assign n31190 = ~n31068 & ~n31083;
  assign n31191 = n75 & n24599;
  assign n31192 = n3020 & n22323;
  assign n31193 = n3023 & n22329;
  assign n31194 = n3028 & n22326;
  assign n31195 = ~n31193 & ~n31194;
  assign n31196 = ~n31192 & n31195;
  assign n31197 = ~n31191 & n31196;
  assign n31198 = ~n13719 & ~n28208;
  assign n31199 =  a[17]  & ~n31198;
  assign n31200 = ~ a[17]  & n31198;
  assign n31201 = ~n31199 & ~n31200;
  assign n31202 = n1143 & n24041;
  assign n31203 = n2719 & n31202;
  assign n31204 = n4785 & n31203;
  assign n31205 = n3282 & n31204;
  assign n31206 = n12924 & n31205;
  assign n31207 = n882 & n31206;
  assign n31208 = n448 & n31207;
  assign n31209 = n279 & n31208;
  assign n31210 = ~n229 & n31209;
  assign n31211 = ~n335 & n31210;
  assign n31212 = ~n299 & n31211;
  assign n31213 = ~n525 & n31212;
  assign n31214 = ~n771 & n31213;
  assign n31215 = n31052 & n31214;
  assign n31216 = ~n31052 & ~n31214;
  assign n31217 = ~n31215 & ~n31216;
  assign n31218 = n31201 & n31217;
  assign n31219 = ~n31201 & ~n31217;
  assign n31220 = ~n31218 & ~n31219;
  assign n31221 = ~n31197 & n31220;
  assign n31222 = n31220 & ~n31221;
  assign n31223 = ~n31197 & ~n31221;
  assign n31224 = ~n31222 & ~n31223;
  assign n31225 = ~n31058 & ~n31224;
  assign n31226 = ~n31224 & ~n31225;
  assign n31227 = ~n31058 & ~n31225;
  assign n31228 = ~n31226 & ~n31227;
  assign n31229 = ~n31190 & ~n31228;
  assign n31230 = ~n31190 & ~n31229;
  assign n31231 = ~n31228 & ~n31229;
  assign n31232 = ~n31230 & ~n31231;
  assign n31233 = n3457 & n22315;
  assign n31234 = n3542 & n22320;
  assign n31235 = n3606 & n22312;
  assign n31236 = ~n31234 & ~n31235;
  assign n31237 = ~n31233 & n31236;
  assign n31238 = n3368 & n25294;
  assign n31239 = n31237 & ~n31238;
  assign n31240 =  a[29]  & ~n31239;
  assign n31241 =  a[29]  & ~n31240;
  assign n31242 = ~n31239 & ~n31240;
  assign n31243 = ~n31241 & ~n31242;
  assign n31244 = ~n31232 & ~n31243;
  assign n31245 = ~n31232 & ~n31244;
  assign n31246 = ~n31243 & ~n31244;
  assign n31247 = ~n31245 & ~n31246;
  assign n31248 = ~n31189 & n31247;
  assign n31249 = n31189 & ~n31247;
  assign n31250 = ~n31248 & ~n31249;
  assign n31251 = n4694 & n27173;
  assign n31252 = n4533 & n26060;
  assign n31253 = n4604 & n26890;
  assign n31254 = ~n31252 & ~n31253;
  assign n31255 = ~n31251 & n31254;
  assign n31256 = n4536 & n27185;
  assign n31257 = n31255 & ~n31256;
  assign n31258 =  a[23]  & ~n31257;
  assign n31259 =  a[23]  & ~n31258;
  assign n31260 = ~n31257 & ~n31258;
  assign n31261 = ~n31259 & ~n31260;
  assign n31262 = ~n31250 & ~n31261;
  assign n31263 = n31250 & n31261;
  assign n31264 = ~n31262 & ~n31263;
  assign n31265 = n31173 & ~n31264;
  assign n31266 = ~n31173 & n31264;
  assign n31267 = ~n31265 & ~n31266;
  assign n31268 = ~n31125 & ~n31138;
  assign n31269 = n5496 & n27964;
  assign n31270 = n4935 & n27442;
  assign n31271 = n5407 & n27698;
  assign n31272 = ~n31270 & ~n31271;
  assign n31273 = ~n31269 & n31272;
  assign n31274 = n4938 & n27976;
  assign n31275 = n31273 & ~n31274;
  assign n31276 =  a[20]  & ~n31275;
  assign n31277 =  a[20]  & ~n31276;
  assign n31278 = ~n31275 & ~n31276;
  assign n31279 = ~n31277 & ~n31278;
  assign n31280 = ~n31268 & ~n31279;
  assign n31281 = ~n31268 & ~n31280;
  assign n31282 = ~n31279 & ~n31280;
  assign n31283 = ~n31281 & ~n31282;
  assign n31284 = ~n31267 & n31283;
  assign n31285 = n31267 & ~n31283;
  assign n31286 = ~n31284 & ~n31285;
  assign n31287 = ~n31172 & n31286;
  assign n31288 = n31172 & ~n31286;
  assign n31289 = ~n31287 & ~n31288;
  assign n31290 = ~n31171 & n31289;
  assign n31291 = n31171 & ~n31289;
  assign n31292 = ~n31290 & ~n31291;
  assign n31293 = ~n31168 & ~n31292;
  assign n31294 = n31168 & n31292;
  assign  result[22]  = ~n31293 & ~n31294;
  assign n31296 = ~n31229 & ~n31244;
  assign n31297 = n75 & ~n25270;
  assign n31298 = n3020 & n22320;
  assign n31299 = n3023 & n22326;
  assign n31300 = n3028 & n22323;
  assign n31301 = ~n31299 & ~n31300;
  assign n31302 = ~n31298 & n31301;
  assign n31303 = ~n31297 & n31302;
  assign n31304 = ~n31216 & ~n31218;
  assign n31305 = n632 & n13014;
  assign n31306 = n2656 & n31305;
  assign n31307 = n6514 & n31306;
  assign n31308 = n2543 & n31307;
  assign n31309 = n3497 & n31308;
  assign n31310 = n29550 & n31309;
  assign n31311 = n423 & n31310;
  assign n31312 = n418 & n31311;
  assign n31313 = n4101 & n31312;
  assign n31314 = ~n330 & n31313;
  assign n31315 = ~n329 & n31314;
  assign n31316 = ~n280 & n31315;
  assign n31317 = ~n203 & n31316;
  assign n31318 = ~n619 & n31317;
  assign n31319 = ~n536 & n31318;
  assign n31320 = ~n31304 & n31319;
  assign n31321 = n31304 & ~n31319;
  assign n31322 = ~n31320 & ~n31321;
  assign n31323 = ~n31303 & n31322;
  assign n31324 = ~n31303 & ~n31323;
  assign n31325 = n31322 & ~n31323;
  assign n31326 = ~n31324 & ~n31325;
  assign n31327 = ~n31221 & ~n31225;
  assign n31328 = n31326 & n31327;
  assign n31329 = ~n31326 & ~n31327;
  assign n31330 = ~n31328 & ~n31329;
  assign n31331 = n3457 & n22309;
  assign n31332 = n3542 & n22312;
  assign n31333 = n3606 & n22315;
  assign n31334 = ~n31332 & ~n31333;
  assign n31335 = ~n31331 & n31334;
  assign n31336 = ~n3368 & n31335;
  assign n31337 = n22529 & n31335;
  assign n31338 = ~n31336 & ~n31337;
  assign n31339 =  a[29]  & ~n31338;
  assign n31340 = ~ a[29]  & n31338;
  assign n31341 = ~n31339 & ~n31340;
  assign n31342 = n31330 & ~n31341;
  assign n31343 = ~n31330 & n31341;
  assign n31344 = ~n31342 & ~n31343;
  assign n31345 = ~n31296 & n31344;
  assign n31346 = n31296 & ~n31344;
  assign n31347 = ~n31345 & ~n31346;
  assign n31348 = n3884 & n26060;
  assign n31349 = n3967 & n26063;
  assign n31350 = n4046 & n26066;
  assign n31351 = ~n31349 & ~n31350;
  assign n31352 = ~n31348 & n31351;
  assign n31353 = n4050 & ~n26088;
  assign n31354 = n31352 & ~n31353;
  assign n31355 =  a[26]  & ~n31354;
  assign n31356 =  a[26]  & ~n31355;
  assign n31357 = ~n31354 & ~n31355;
  assign n31358 = ~n31356 & ~n31357;
  assign n31359 = n31347 & ~n31358;
  assign n31360 = n31347 & ~n31359;
  assign n31361 = ~n31358 & ~n31359;
  assign n31362 = ~n31360 & ~n31361;
  assign n31363 = ~n31189 & ~n31247;
  assign n31364 = ~n31186 & ~n31363;
  assign n31365 = ~n31362 & ~n31364;
  assign n31366 = ~n31362 & ~n31365;
  assign n31367 = ~n31364 & ~n31365;
  assign n31368 = ~n31366 & ~n31367;
  assign n31369 = n4694 & n27442;
  assign n31370 = n4533 & n26890;
  assign n31371 = n4604 & n27173;
  assign n31372 = ~n31370 & ~n31371;
  assign n31373 = ~n31369 & n31372;
  assign n31374 = n4536 & n27455;
  assign n31375 = n31373 & ~n31374;
  assign n31376 =  a[23]  & ~n31375;
  assign n31377 =  a[23]  & ~n31376;
  assign n31378 = ~n31375 & ~n31376;
  assign n31379 = ~n31377 & ~n31378;
  assign n31380 = ~n31368 & ~n31379;
  assign n31381 = ~n31368 & ~n31380;
  assign n31382 = ~n31379 & ~n31380;
  assign n31383 = ~n31381 & ~n31382;
  assign n31384 = ~n31262 & ~n31266;
  assign n31385 = n31383 & n31384;
  assign n31386 = ~n31383 & ~n31384;
  assign n31387 = ~n31385 & ~n31386;
  assign n31388 = n5496 & ~n28208;
  assign n31389 = n4935 & n27698;
  assign n31390 = n5407 & n27964;
  assign n31391 = ~n31389 & ~n31390;
  assign n31392 = ~n31388 & n31391;
  assign n31393 = n4938 & ~n28223;
  assign n31394 = n31392 & ~n31393;
  assign n31395 =  a[20]  & ~n31394;
  assign n31396 =  a[20]  & ~n31395;
  assign n31397 = ~n31394 & ~n31395;
  assign n31398 = ~n31396 & ~n31397;
  assign n31399 = n31387 & ~n31398;
  assign n31400 = n31387 & ~n31399;
  assign n31401 = ~n31398 & ~n31399;
  assign n31402 = ~n31400 & ~n31401;
  assign n31403 = ~n31280 & ~n31285;
  assign n31404 = ~n31402 & ~n31403;
  assign n31405 = ~n31402 & ~n31404;
  assign n31406 = ~n31403 & ~n31404;
  assign n31407 = ~n31405 & ~n31406;
  assign n31408 = ~n31287 & ~n31290;
  assign n31409 = n31407 & n31408;
  assign n31410 = ~n31407 & ~n31408;
  assign n31411 = ~n31409 & ~n31410;
  assign n31412 = ~n31294 & n31411;
  assign n31413 = n31294 & ~n31411;
  assign  result[23]  = n31412 | n31413;
  assign n31415 = n31294 & n31411;
  assign n31416 = n75 & ~n25315;
  assign n31417 = n3020 & n22312;
  assign n31418 = n3023 & n22323;
  assign n31419 = n3028 & n22320;
  assign n31420 = ~n31418 & ~n31419;
  assign n31421 = ~n31417 & n31420;
  assign n31422 = ~n31416 & n31421;
  assign n31423 = n12941 & n31036;
  assign n31424 = n4366 & n31423;
  assign n31425 = n6561 & n31424;
  assign n31426 = n3259 & n31425;
  assign n31427 = n2651 & n31426;
  assign n31428 = n2683 & n31427;
  assign n31429 = n230 & n31428;
  assign n31430 = n488 & n31429;
  assign n31431 = n28688 & n31430;
  assign n31432 = ~n602 & n31431;
  assign n31433 = ~n1101 & n31432;
  assign n31434 = ~n142 & n31433;
  assign n31435 = ~n125 & n31434;
  assign n31436 = ~n31319 & n31435;
  assign n31437 = n31319 & ~n31435;
  assign n31438 = ~n31422 & ~n31437;
  assign n31439 = ~n31436 & n31438;
  assign n31440 = ~n31422 & ~n31439;
  assign n31441 = ~n31437 & ~n31439;
  assign n31442 = ~n31436 & n31441;
  assign n31443 = ~n31440 & ~n31442;
  assign n31444 = ~n31320 & ~n31323;
  assign n31445 = n31443 & n31444;
  assign n31446 = ~n31443 & ~n31444;
  assign n31447 = ~n31445 & ~n31446;
  assign n31448 = ~n31329 & ~n31342;
  assign n31449 = ~n31447 & n31448;
  assign n31450 = n31447 & ~n31448;
  assign n31451 = ~n31449 & ~n31450;
  assign n31452 = n3457 & n26063;
  assign n31453 = n3542 & n22315;
  assign n31454 = n3606 & n22309;
  assign n31455 = ~n31453 & ~n31454;
  assign n31456 = ~n31452 & n31455;
  assign n31457 = n3368 & ~n26604;
  assign n31458 = n31456 & ~n31457;
  assign n31459 =  a[29]  & ~n31458;
  assign n31460 =  a[29]  & ~n31459;
  assign n31461 = ~n31458 & ~n31459;
  assign n31462 = ~n31460 & ~n31461;
  assign n31463 = n31451 & ~n31462;
  assign n31464 = n31451 & ~n31463;
  assign n31465 = ~n31462 & ~n31463;
  assign n31466 = ~n31464 & ~n31465;
  assign n31467 = n3884 & n26890;
  assign n31468 = n3967 & n26066;
  assign n31469 = n4046 & n26060;
  assign n31470 = ~n31468 & ~n31469;
  assign n31471 = ~n31467 & n31470;
  assign n31472 = n4050 & ~n26904;
  assign n31473 = n31471 & ~n31472;
  assign n31474 =  a[26]  & ~n31473;
  assign n31475 =  a[26]  & ~n31474;
  assign n31476 = ~n31473 & ~n31474;
  assign n31477 = ~n31475 & ~n31476;
  assign n31478 = ~n31466 & ~n31477;
  assign n31479 = ~n31466 & ~n31478;
  assign n31480 = ~n31477 & ~n31478;
  assign n31481 = ~n31479 & ~n31480;
  assign n31482 = ~n31345 & ~n31359;
  assign n31483 = n31481 & n31482;
  assign n31484 = ~n31481 & ~n31482;
  assign n31485 = ~n31483 & ~n31484;
  assign n31486 = n4694 & n27698;
  assign n31487 = n4533 & n27173;
  assign n31488 = n4604 & n27442;
  assign n31489 = ~n31487 & ~n31488;
  assign n31490 = ~n31486 & n31489;
  assign n31491 = n4536 & ~n27713;
  assign n31492 = n31490 & ~n31491;
  assign n31493 =  a[23]  & ~n31492;
  assign n31494 =  a[23]  & ~n31493;
  assign n31495 = ~n31492 & ~n31493;
  assign n31496 = ~n31494 & ~n31495;
  assign n31497 = n31485 & ~n31496;
  assign n31498 = n31485 & ~n31497;
  assign n31499 = ~n31496 & ~n31497;
  assign n31500 = ~n31498 & ~n31499;
  assign n31501 = ~n31365 & ~n31380;
  assign n31502 = ~n13439 & ~n28208;
  assign n31503 = n4935 & n27964;
  assign n31504 = ~n31502 & ~n31503;
  assign n31505 = ~n4938 & n31504;
  assign n31506 = n28221 & n31504;
  assign n31507 = ~n31505 & ~n31506;
  assign n31508 =  a[20]  & ~n31507;
  assign n31509 = ~ a[20]  & n31507;
  assign n31510 = ~n31508 & ~n31509;
  assign n31511 = ~n31501 & ~n31510;
  assign n31512 = n31501 & n31510;
  assign n31513 = ~n31511 & ~n31512;
  assign n31514 = ~n31500 & n31513;
  assign n31515 = ~n31500 & ~n31514;
  assign n31516 = n31513 & ~n31514;
  assign n31517 = ~n31515 & ~n31516;
  assign n31518 = ~n31386 & ~n31399;
  assign n31519 = n31517 & n31518;
  assign n31520 = ~n31517 & ~n31518;
  assign n31521 = ~n31519 & ~n31520;
  assign n31522 = ~n31404 & ~n31410;
  assign n31523 = ~n31521 & n31522;
  assign n31524 = n31521 & ~n31522;
  assign n31525 = ~n31523 & ~n31524;
  assign n31526 = n31415 & n31525;
  assign n31527 = ~n31415 & ~n31525;
  assign  result[24]  = ~n31526 & ~n31527;
  assign n31529 = ~n31520 & ~n31524;
  assign n31530 = ~n31511 & ~n31514;
  assign n31531 = n75 & n25294;
  assign n31532 = n3020 & n22315;
  assign n31533 = n3023 & n22320;
  assign n31534 = n3028 & n22312;
  assign n31535 = ~n31533 & ~n31534;
  assign n31536 = ~n31532 & n31535;
  assign n31537 = ~n31531 & n31536;
  assign n31538 = ~n13441 & ~n28208;
  assign n31539 =  a[20]  & ~n31538;
  assign n31540 = ~ a[20]  & n31538;
  assign n31541 = ~n31539 & ~n31540;
  assign n31542 = n2753 & n3370;
  assign n31543 = n530 & n31542;
  assign n31544 = n15050 & n31543;
  assign n31545 = n15953 & n31544;
  assign n31546 = n4293 & n31545;
  assign n31547 = n1008 & n31546;
  assign n31548 = n805 & n31547;
  assign n31549 = n539 & n31548;
  assign n31550 = n2506 & n31549;
  assign n31551 = n615 & n31550;
  assign n31552 = n1574 & n31551;
  assign n31553 = ~n558 & n31552;
  assign n31554 = ~n420 & n31553;
  assign n31555 = ~n189 & n31554;
  assign n31556 = ~n716 & n31555;
  assign n31557 = ~n452 & n31556;
  assign n31558 = ~n201 & n31557;
  assign n31559 = n31319 & n31558;
  assign n31560 = ~n31319 & ~n31558;
  assign n31561 = ~n31559 & ~n31560;
  assign n31562 = n31541 & n31561;
  assign n31563 = ~n31541 & ~n31561;
  assign n31564 = ~n31562 & ~n31563;
  assign n31565 = ~n31441 & n31564;
  assign n31566 = n31441 & ~n31564;
  assign n31567 = ~n31565 & ~n31566;
  assign n31568 = ~n31537 & n31567;
  assign n31569 = n31567 & ~n31568;
  assign n31570 = ~n31537 & ~n31568;
  assign n31571 = ~n31569 & ~n31570;
  assign n31572 = ~n31446 & ~n31450;
  assign n31573 = n31571 & n31572;
  assign n31574 = ~n31571 & ~n31572;
  assign n31575 = ~n31573 & ~n31574;
  assign n31576 = n3457 & n26066;
  assign n31577 = n3542 & n22309;
  assign n31578 = n3606 & n26063;
  assign n31579 = ~n31577 & ~n31578;
  assign n31580 = ~n31576 & n31579;
  assign n31581 = n3368 & ~n26624;
  assign n31582 = n31580 & ~n31581;
  assign n31583 =  a[29]  & ~n31582;
  assign n31584 =  a[29]  & ~n31583;
  assign n31585 = ~n31582 & ~n31583;
  assign n31586 = ~n31584 & ~n31585;
  assign n31587 = n31575 & ~n31586;
  assign n31588 = n31575 & ~n31587;
  assign n31589 = ~n31586 & ~n31587;
  assign n31590 = ~n31588 & ~n31589;
  assign n31591 = n3884 & n27173;
  assign n31592 = n3967 & n26060;
  assign n31593 = n4046 & n26890;
  assign n31594 = ~n31592 & ~n31593;
  assign n31595 = ~n31591 & n31594;
  assign n31596 = n4050 & n27185;
  assign n31597 = n31595 & ~n31596;
  assign n31598 =  a[26]  & ~n31597;
  assign n31599 =  a[26]  & ~n31598;
  assign n31600 = ~n31597 & ~n31598;
  assign n31601 = ~n31599 & ~n31600;
  assign n31602 = ~n31590 & ~n31601;
  assign n31603 = ~n31590 & ~n31602;
  assign n31604 = ~n31601 & ~n31602;
  assign n31605 = ~n31603 & ~n31604;
  assign n31606 = ~n31463 & ~n31478;
  assign n31607 = n31605 & n31606;
  assign n31608 = ~n31605 & ~n31606;
  assign n31609 = ~n31607 & ~n31608;
  assign n31610 = ~n31484 & ~n31497;
  assign n31611 = n4694 & n27964;
  assign n31612 = n4533 & n27442;
  assign n31613 = n4604 & n27698;
  assign n31614 = ~n31612 & ~n31613;
  assign n31615 = ~n31611 & n31614;
  assign n31616 = n4536 & n27976;
  assign n31617 = n31615 & ~n31616;
  assign n31618 =  a[23]  & ~n31617;
  assign n31619 =  a[23]  & ~n31618;
  assign n31620 = ~n31617 & ~n31618;
  assign n31621 = ~n31619 & ~n31620;
  assign n31622 = ~n31610 & ~n31621;
  assign n31623 = ~n31610 & ~n31622;
  assign n31624 = ~n31621 & ~n31622;
  assign n31625 = ~n31623 & ~n31624;
  assign n31626 = ~n31609 & n31625;
  assign n31627 = n31609 & ~n31625;
  assign n31628 = ~n31626 & ~n31627;
  assign n31629 = ~n31530 & n31628;
  assign n31630 = n31530 & ~n31628;
  assign n31631 = ~n31629 & ~n31630;
  assign n31632 = ~n31529 & n31631;
  assign n31633 = n31529 & ~n31631;
  assign n31634 = ~n31632 & ~n31633;
  assign n31635 = ~n31526 & ~n31634;
  assign n31636 = n31526 & n31634;
  assign  result[25]  = ~n31635 & ~n31636;
  assign n31638 = ~n31574 & ~n31587;
  assign n31639 = n75 & ~n22529;
  assign n31640 = n3020 & n22309;
  assign n31641 = n3023 & n22312;
  assign n31642 = n3028 & n22315;
  assign n31643 = ~n31641 & ~n31642;
  assign n31644 = ~n31640 & n31643;
  assign n31645 = ~n31639 & n31644;
  assign n31646 = ~n31560 & ~n31562;
  assign n31647 = n1740 & n4828;
  assign n31648 = n1604 & n31647;
  assign n31649 = n1640 & n31648;
  assign n31650 = n14534 & n31649;
  assign n31651 = n1029 & n31650;
  assign n31652 = n3282 & n31651;
  assign n31653 = n1679 & n31652;
  assign n31654 = n3039 & n31653;
  assign n31655 = n16055 & n31654;
  assign n31656 = n1252 & n31655;
  assign n31657 = ~n1246 & n31656;
  assign n31658 = ~n602 & n31657;
  assign n31659 = ~n145 & n31658;
  assign n31660 = ~n298 & n31659;
  assign n31661 = ~n222 & n31660;
  assign n31662 = ~n31646 & n31661;
  assign n31663 = n31646 & ~n31661;
  assign n31664 = ~n31662 & ~n31663;
  assign n31665 = ~n31645 & n31664;
  assign n31666 = ~n31645 & ~n31665;
  assign n31667 = n31664 & ~n31665;
  assign n31668 = ~n31666 & ~n31667;
  assign n31669 = ~n31565 & ~n31568;
  assign n31670 = n31668 & n31669;
  assign n31671 = ~n31668 & ~n31669;
  assign n31672 = ~n31670 & ~n31671;
  assign n31673 = n3457 & n26060;
  assign n31674 = n3542 & n26063;
  assign n31675 = n3606 & n26066;
  assign n31676 = ~n31674 & ~n31675;
  assign n31677 = ~n31673 & n31676;
  assign n31678 = ~n3368 & n31677;
  assign n31679 = n26088 & n31677;
  assign n31680 = ~n31678 & ~n31679;
  assign n31681 =  a[29]  & ~n31680;
  assign n31682 = ~ a[29]  & n31680;
  assign n31683 = ~n31681 & ~n31682;
  assign n31684 = n31672 & ~n31683;
  assign n31685 = ~n31672 & n31683;
  assign n31686 = ~n31684 & ~n31685;
  assign n31687 = ~n31638 & n31686;
  assign n31688 = n31638 & ~n31686;
  assign n31689 = ~n31687 & ~n31688;
  assign n31690 = n3884 & n27442;
  assign n31691 = n3967 & n26890;
  assign n31692 = n4046 & n27173;
  assign n31693 = ~n31691 & ~n31692;
  assign n31694 = ~n31690 & n31693;
  assign n31695 = n4050 & n27455;
  assign n31696 = n31694 & ~n31695;
  assign n31697 =  a[26]  & ~n31696;
  assign n31698 =  a[26]  & ~n31697;
  assign n31699 = ~n31696 & ~n31697;
  assign n31700 = ~n31698 & ~n31699;
  assign n31701 = n31689 & ~n31700;
  assign n31702 = n31689 & ~n31701;
  assign n31703 = ~n31700 & ~n31701;
  assign n31704 = ~n31702 & ~n31703;
  assign n31705 = ~n31602 & ~n31608;
  assign n31706 = n31704 & n31705;
  assign n31707 = ~n31704 & ~n31705;
  assign n31708 = ~n31706 & ~n31707;
  assign n31709 = n4694 & ~n28208;
  assign n31710 = n4533 & n27698;
  assign n31711 = n4604 & n27964;
  assign n31712 = ~n31710 & ~n31711;
  assign n31713 = ~n31709 & n31712;
  assign n31714 = n4536 & ~n28223;
  assign n31715 = n31713 & ~n31714;
  assign n31716 =  a[23]  & ~n31715;
  assign n31717 =  a[23]  & ~n31716;
  assign n31718 = ~n31715 & ~n31716;
  assign n31719 = ~n31717 & ~n31718;
  assign n31720 = n31708 & ~n31719;
  assign n31721 = n31708 & ~n31720;
  assign n31722 = ~n31719 & ~n31720;
  assign n31723 = ~n31721 & ~n31722;
  assign n31724 = ~n31622 & ~n31627;
  assign n31725 = ~n31723 & ~n31724;
  assign n31726 = ~n31723 & ~n31725;
  assign n31727 = ~n31724 & ~n31725;
  assign n31728 = ~n31726 & ~n31727;
  assign n31729 = ~n31629 & ~n31632;
  assign n31730 = n31728 & n31729;
  assign n31731 = ~n31728 & ~n31729;
  assign n31732 = ~n31730 & ~n31731;
  assign n31733 = n31636 & ~n31732;
  assign n31734 = ~n31636 & n31732;
  assign  result[26]  = n31733 | n31734;
  assign n31736 = ~n31662 & ~n31665;
  assign n31737 = n3459 & n13016;
  assign n31738 = n1070 & n31737;
  assign n31739 = n15882 & n31738;
  assign n31740 = n25863 & n31739;
  assign n31741 = n4232 & n31740;
  assign n31742 = n2651 & n31741;
  assign n31743 = n29538 & n31742;
  assign n31744 = n285 & n31743;
  assign n31745 = n1252 & n31744;
  assign n31746 = n720 & n31745;
  assign n31747 = n22762 & n31746;
  assign n31748 = ~n334 & n31747;
  assign n31749 = ~n233 & n31748;
  assign n31750 = ~n302 & n31749;
  assign n31751 = ~n714 & n31750;
  assign n31752 = n31661 & ~n31751;
  assign n31753 = ~n31661 & n31751;
  assign n31754 = ~n31736 & ~n31753;
  assign n31755 = ~n31752 & n31754;
  assign n31756 = ~n31736 & ~n31755;
  assign n31757 = ~n31753 & ~n31755;
  assign n31758 = ~n31752 & n31757;
  assign n31759 = ~n31756 & ~n31758;
  assign n31760 = n75 & ~n26604;
  assign n31761 = n3020 & n26063;
  assign n31762 = n3023 & n22315;
  assign n31763 = n3028 & n22309;
  assign n31764 = ~n31762 & ~n31763;
  assign n31765 = ~n31761 & n31764;
  assign n31766 = ~n31760 & n31765;
  assign n31767 = ~n31759 & ~n31766;
  assign n31768 = ~n31759 & ~n31767;
  assign n31769 = ~n31766 & ~n31767;
  assign n31770 = ~n31768 & ~n31769;
  assign n31771 = ~n31671 & ~n31684;
  assign n31772 = n31770 & n31771;
  assign n31773 = ~n31770 & ~n31771;
  assign n31774 = ~n31772 & ~n31773;
  assign n31775 = n3457 & n26890;
  assign n31776 = n3542 & n26066;
  assign n31777 = n3606 & n26060;
  assign n31778 = ~n31776 & ~n31777;
  assign n31779 = ~n31775 & n31778;
  assign n31780 = n3368 & ~n26904;
  assign n31781 = n31779 & ~n31780;
  assign n31782 =  a[29]  & ~n31781;
  assign n31783 =  a[29]  & ~n31782;
  assign n31784 = ~n31781 & ~n31782;
  assign n31785 = ~n31783 & ~n31784;
  assign n31786 = n31774 & ~n31785;
  assign n31787 = n31774 & ~n31786;
  assign n31788 = ~n31785 & ~n31786;
  assign n31789 = ~n31787 & ~n31788;
  assign n31790 = n3884 & n27698;
  assign n31791 = n3967 & n27173;
  assign n31792 = n4046 & n27442;
  assign n31793 = ~n31791 & ~n31792;
  assign n31794 = ~n31790 & n31793;
  assign n31795 = n4050 & ~n27713;
  assign n31796 = n31794 & ~n31795;
  assign n31797 =  a[26]  & ~n31796;
  assign n31798 =  a[26]  & ~n31797;
  assign n31799 = ~n31796 & ~n31797;
  assign n31800 = ~n31798 & ~n31799;
  assign n31801 = ~n31789 & ~n31800;
  assign n31802 = ~n31789 & ~n31801;
  assign n31803 = ~n31800 & ~n31801;
  assign n31804 = ~n31802 & ~n31803;
  assign n31805 = ~n31687 & ~n31701;
  assign n31806 = ~n13938 & ~n28208;
  assign n31807 = n4533 & n27964;
  assign n31808 = ~n31806 & ~n31807;
  assign n31809 = ~n4536 & n31808;
  assign n31810 = n28221 & n31808;
  assign n31811 = ~n31809 & ~n31810;
  assign n31812 =  a[23]  & ~n31811;
  assign n31813 = ~ a[23]  & n31811;
  assign n31814 = ~n31812 & ~n31813;
  assign n31815 = ~n31805 & ~n31814;
  assign n31816 = n31805 & n31814;
  assign n31817 = ~n31815 & ~n31816;
  assign n31818 = ~n31804 & n31817;
  assign n31819 = ~n31804 & ~n31818;
  assign n31820 = n31817 & ~n31818;
  assign n31821 = ~n31819 & ~n31820;
  assign n31822 = ~n31707 & ~n31720;
  assign n31823 = n31821 & n31822;
  assign n31824 = ~n31821 & ~n31822;
  assign n31825 = ~n31823 & ~n31824;
  assign n31826 = ~n31725 & ~n31731;
  assign n31827 = ~n31825 & n31826;
  assign n31828 = n31825 & ~n31826;
  assign n31829 = ~n31827 & ~n31828;
  assign n31830 = n31636 & n31732;
  assign n31831 = n31829 & n31830;
  assign n31832 = ~n31829 & ~n31830;
  assign  result[27]  = ~n31831 & ~n31832;
  assign n31834 = ~n31824 & ~n31828;
  assign n31835 = ~n31815 & ~n31818;
  assign n31836 = ~n31786 & ~n31801;
  assign n31837 = n3884 & n27964;
  assign n31838 = n3967 & n27442;
  assign n31839 = n4046 & n27698;
  assign n31840 = ~n31838 & ~n31839;
  assign n31841 = ~n31837 & n31840;
  assign n31842 = n4050 & n27976;
  assign n31843 = n31841 & ~n31842;
  assign n31844 =  a[26]  & ~n31843;
  assign n31845 =  a[26]  & ~n31844;
  assign n31846 = ~n31843 & ~n31844;
  assign n31847 = ~n31845 & ~n31846;
  assign n31848 = ~n31836 & ~n31847;
  assign n31849 = ~n31836 & ~n31848;
  assign n31850 = ~n31847 & ~n31848;
  assign n31851 = ~n31849 & ~n31850;
  assign n31852 = n75 & ~n26624;
  assign n31853 = n3020 & n26066;
  assign n31854 = n3023 & n22309;
  assign n31855 = n3028 & n26063;
  assign n31856 = ~n31854 & ~n31855;
  assign n31857 = ~n31853 & n31856;
  assign n31858 = ~n31852 & n31857;
  assign n31859 = ~n22248 & ~n28208;
  assign n31860 =  a[23]  & ~n31859;
  assign n31861 = ~ a[23]  & n31859;
  assign n31862 = ~n31860 & ~n31861;
  assign n31863 = n4799 & n13161;
  assign n31864 = n1155 & n31863;
  assign n31865 = n4003 & n31864;
  assign n31866 = n3866 & n31865;
  assign n31867 = n288 & n31866;
  assign n31868 = n937 & n31867;
  assign n31869 = n1478 & n31868;
  assign n31870 = n193 & n31869;
  assign n31871 = ~n509 & n31870;
  assign n31872 = ~n1011 & n31871;
  assign n31873 = ~n228 & n31872;
  assign n31874 = ~n825 & n31873;
  assign n31875 = ~n568 & n31874;
  assign n31876 = ~n519 & n31875;
  assign n31877 = n31751 & n31876;
  assign n31878 = ~n31751 & ~n31876;
  assign n31879 = ~n31877 & ~n31878;
  assign n31880 = n31862 & n31879;
  assign n31881 = ~n31862 & ~n31879;
  assign n31882 = ~n31880 & ~n31881;
  assign n31883 = ~n31757 & n31882;
  assign n31884 = n31757 & ~n31882;
  assign n31885 = ~n31883 & ~n31884;
  assign n31886 = ~n31858 & n31885;
  assign n31887 = n31885 & ~n31886;
  assign n31888 = ~n31858 & ~n31886;
  assign n31889 = ~n31887 & ~n31888;
  assign n31890 = ~n31767 & ~n31773;
  assign n31891 = n31889 & n31890;
  assign n31892 = ~n31889 & ~n31890;
  assign n31893 = ~n31891 & ~n31892;
  assign n31894 = n3457 & n27173;
  assign n31895 = n3542 & n26060;
  assign n31896 = n3606 & n26890;
  assign n31897 = ~n31895 & ~n31896;
  assign n31898 = ~n31894 & n31897;
  assign n31899 = n3368 & n27185;
  assign n31900 = n31898 & ~n31899;
  assign n31901 =  a[29]  & ~n31900;
  assign n31902 =  a[29]  & ~n31901;
  assign n31903 = ~n31900 & ~n31901;
  assign n31904 = ~n31902 & ~n31903;
  assign n31905 = n31893 & ~n31904;
  assign n31906 = n31893 & ~n31905;
  assign n31907 = ~n31904 & ~n31905;
  assign n31908 = ~n31906 & ~n31907;
  assign n31909 = ~n31851 & n31908;
  assign n31910 = n31851 & ~n31908;
  assign n31911 = ~n31909 & ~n31910;
  assign n31912 = ~n31835 & ~n31911;
  assign n31913 = n31835 & n31911;
  assign n31914 = ~n31912 & ~n31913;
  assign n31915 = ~n31834 & n31914;
  assign n31916 = n31834 & ~n31914;
  assign n31917 = ~n31915 & ~n31916;
  assign n31918 = ~n31831 & ~n31917;
  assign n31919 = n31831 & n31917;
  assign  result[28]  = ~n31918 & ~n31919;
  assign n31921 = ~n31892 & ~n31905;
  assign n31922 = n75 & ~n26088;
  assign n31923 = n3020 & n26060;
  assign n31924 = n3023 & n26063;
  assign n31925 = n3028 & n26066;
  assign n31926 = ~n31924 & ~n31925;
  assign n31927 = ~n31923 & n31926;
  assign n31928 = ~n31922 & n31927;
  assign n31929 = ~n31878 & ~n31880;
  assign n31930 = n1738 & n15012;
  assign n31931 = n3438 & n31930;
  assign n31932 = n6610 & n31931;
  assign n31933 = n26016 & n31932;
  assign n31934 = n15880 & n31933;
  assign n31935 = n3939 & n31934;
  assign n31936 = n3997 & n31935;
  assign n31937 = n1183 & n31936;
  assign n31938 = n1531 & n31937;
  assign n31939 = n1366 & n31938;
  assign n31940 = n1783 & n31939;
  assign n31941 = n100 & n31940;
  assign n31942 = ~n420 & n31941;
  assign n31943 = ~n466 & n31942;
  assign n31944 = ~n298 & n31943;
  assign n31945 = ~n251 & n31944;
  assign n31946 = ~n31929 & n31945;
  assign n31947 = n31929 & ~n31945;
  assign n31948 = ~n31946 & ~n31947;
  assign n31949 = ~n31928 & n31948;
  assign n31950 = ~n31928 & ~n31949;
  assign n31951 = n31948 & ~n31949;
  assign n31952 = ~n31950 & ~n31951;
  assign n31953 = ~n31883 & ~n31886;
  assign n31954 = n31952 & n31953;
  assign n31955 = ~n31952 & ~n31953;
  assign n31956 = ~n31954 & ~n31955;
  assign n31957 = n3457 & n27442;
  assign n31958 = n3542 & n26890;
  assign n31959 = n3606 & n27173;
  assign n31960 = ~n31958 & ~n31959;
  assign n31961 = ~n31957 & n31960;
  assign n31962 = ~n3368 & n31961;
  assign n31963 = ~n27455 & n31961;
  assign n31964 = ~n31962 & ~n31963;
  assign n31965 =  a[29]  & ~n31964;
  assign n31966 = ~ a[29]  & n31964;
  assign n31967 = ~n31965 & ~n31966;
  assign n31968 = n31956 & ~n31967;
  assign n31969 = ~n31956 & n31967;
  assign n31970 = ~n31968 & ~n31969;
  assign n31971 = ~n31921 & n31970;
  assign n31972 = n31921 & ~n31970;
  assign n31973 = ~n31971 & ~n31972;
  assign n31974 = n3884 & ~n28208;
  assign n31975 = n3967 & n27698;
  assign n31976 = n4046 & n27964;
  assign n31977 = ~n31975 & ~n31976;
  assign n31978 = ~n31974 & n31977;
  assign n31979 = n4050 & ~n28223;
  assign n31980 = n31978 & ~n31979;
  assign n31981 =  a[26]  & ~n31980;
  assign n31982 =  a[26]  & ~n31981;
  assign n31983 = ~n31980 & ~n31981;
  assign n31984 = ~n31982 & ~n31983;
  assign n31985 = n31973 & ~n31984;
  assign n31986 = n31973 & ~n31985;
  assign n31987 = ~n31984 & ~n31985;
  assign n31988 = ~n31986 & ~n31987;
  assign n31989 = ~n31851 & ~n31908;
  assign n31990 = ~n31848 & ~n31989;
  assign n31991 = ~n31988 & ~n31990;
  assign n31992 = ~n31988 & ~n31991;
  assign n31993 = ~n31990 & ~n31991;
  assign n31994 = ~n31992 & ~n31993;
  assign n31995 = ~n31912 & ~n31915;
  assign n31996 = n31994 & n31995;
  assign n31997 = ~n31994 & ~n31995;
  assign n31998 = ~n31996 & ~n31997;
  assign n31999 = ~n31919 & n31998;
  assign n32000 = n31919 & ~n31998;
  assign  result[29]  = n31999 | n32000;
  assign n32002 = n31919 & n31998;
  assign n32003 = ~n31991 & ~n31997;
  assign n32004 = ~n31971 & ~n31985;
  assign n32005 = ~n31946 & ~n31949;
  assign n32006 = n4009 & n13075;
  assign n32007 = n3848 & n32006;
  assign n32008 = n3839 & n32007;
  assign n32009 = n2273 & n32008;
  assign n32010 = n26016 & n32009;
  assign n32011 = n3984 & n32010;
  assign n32012 = ~n825 & n32011;
  assign n32013 = ~n31945 & n32012;
  assign n32014 = n31945 & ~n32012;
  assign n32015 = ~n32005 & ~n32014;
  assign n32016 = ~n32013 & n32015;
  assign n32017 = ~n32005 & ~n32016;
  assign n32018 = ~n32014 & ~n32016;
  assign n32019 = ~n32013 & n32018;
  assign n32020 = ~n32017 & ~n32019;
  assign n32021 = n75 & ~n26904;
  assign n32022 = n3020 & n26890;
  assign n32023 = n3023 & n26066;
  assign n32024 = n3028 & n26060;
  assign n32025 = ~n32023 & ~n32024;
  assign n32026 = ~n32022 & n32025;
  assign n32027 = ~n32021 & n32026;
  assign n32028 = ~n32020 & ~n32027;
  assign n32029 = ~n32020 & ~n32028;
  assign n32030 = ~n32027 & ~n32028;
  assign n32031 = ~n32029 & ~n32030;
  assign n32032 = ~n31955 & ~n31968;
  assign n32033 = n32031 & n32032;
  assign n32034 = ~n32031 & ~n32032;
  assign n32035 = ~n32033 & ~n32034;
  assign n32036 = ~n25957 & ~n28208;
  assign n32037 = n3967 & n27964;
  assign n32038 = ~n32036 & ~n32037;
  assign n32039 = n4050 & ~n28221;
  assign n32040 = n32038 & ~n32039;
  assign n32041 =  a[26]  & ~n32040;
  assign n32042 = ~n32040 & ~n32041;
  assign n32043 =  a[26]  & ~n32041;
  assign n32044 = ~n32042 & ~n32043;
  assign n32045 = n3457 & n27698;
  assign n32046 = n3542 & n27173;
  assign n32047 = n3606 & n27442;
  assign n32048 = ~n32046 & ~n32047;
  assign n32049 = ~n32045 & n32048;
  assign n32050 = n3368 & ~n27713;
  assign n32051 = n32049 & ~n32050;
  assign n32052 =  a[29]  & ~n32051;
  assign n32053 =  a[29]  & ~n32052;
  assign n32054 = ~n32051 & ~n32052;
  assign n32055 = ~n32053 & ~n32054;
  assign n32056 = ~n32044 & ~n32055;
  assign n32057 = ~n32044 & ~n32056;
  assign n32058 = ~n32055 & ~n32056;
  assign n32059 = ~n32057 & ~n32058;
  assign n32060 = ~n32035 & n32059;
  assign n32061 = n32035 & ~n32059;
  assign n32062 = ~n32060 & ~n32061;
  assign n32063 = ~n32004 & n32062;
  assign n32064 = n32004 & ~n32062;
  assign n32065 = ~n32063 & ~n32064;
  assign n32066 = ~n32003 & n32065;
  assign n32067 = n32003 & ~n32065;
  assign n32068 = ~n32066 & ~n32067;
  assign n32069 = ~n32002 & ~n32068;
  assign n32070 = n32002 & n32068;
  assign  result[30]  = ~n32069 & ~n32070;
  assign n32072 = ~n32063 & ~n32066;
  assign n32073 = n3457 & n27964;
  assign n32074 = n3542 & n27442;
  assign n32075 = n3606 & n27698;
  assign n32076 = ~n32074 & ~n32075;
  assign n32077 = ~n32073 & n32076;
  assign n32078 = n3368 & n27976;
  assign n32079 = n32077 & ~n32078;
  assign n32080 = ~n32028 & ~n32034;
  assign n32081 =  a[29]  & ~n32080;
  assign n32082 = ~ a[29]  & n32080;
  assign n32083 = ~n32081 & ~n32082;
  assign n32084 = n32079 & n32083;
  assign n32085 = ~n32079 & ~n32083;
  assign n32086 = ~n32084 & ~n32085;
  assign n32087 = n75 & n27185;
  assign n32088 = n3020 & n27173;
  assign n32089 = n3023 & n26060;
  assign n32090 = n3028 & n26890;
  assign n32091 = ~n32089 & ~n32090;
  assign n32092 = ~n32088 & n32091;
  assign n32093 = ~n32087 & n32092;
  assign n32094 = n32018 & ~n32093;
  assign n32095 = ~n32018 & n32093;
  assign n32096 = ~n32094 & ~n32095;
  assign n32097 = n32086 & ~n32096;
  assign n32098 = ~n32086 & n32096;
  assign n32099 = ~n32097 & ~n32098;
  assign n32100 = ~n32056 & ~n32061;
  assign n32101 = n3874 & n4511;
  assign n32102 = ~n601 & n32101;
  assign n32103 =  a[26]  & ~n32102;
  assign n32104 = ~ a[26]  & n32102;
  assign n32105 = ~n32103 & ~n32104;
  assign n32106 = ~n26010 & ~n28208;
  assign n32107 = n31945 & ~n32106;
  assign n32108 = ~n31945 & n32106;
  assign n32109 = ~n32107 & ~n32108;
  assign n32110 = n32105 & n32109;
  assign n32111 = ~n32105 & ~n32109;
  assign n32112 = ~n32110 & ~n32111;
  assign n32113 = n32100 & ~n32112;
  assign n32114 = ~n32100 & n32112;
  assign n32115 = ~n32113 & ~n32114;
  assign n32116 = n32099 & n32115;
  assign n32117 = ~n32099 & ~n32115;
  assign n32118 = ~n32116 & ~n32117;
  assign n32119 = ~n32072 & ~n32118;
  assign n32120 = n32072 & n32118;
  assign n32121 = ~n32119 & ~n32120;
  assign n32122 = n32070 & n32121;
  assign n32123 = ~n32070 & ~n32121;
  assign  result[31]  = n32122 | n32123;
endmodule


