module dec ( count , selectp1 , selectp2   );
  input  [7:0] count ;
  output wire [127:0] selectp1, selectp2;
  wire n265, n266, n267, n268, n269, n270, n272, n273, n275, n276, n278,
    n280, n281, n283, n284, n286, n288, n290, n291, n293, n295, n296, n298,
    n300, n302, n304, n306, n308, n309, n326, n327, n344, n345, n362, n363,
    n380, n397, n414, n431, n432, n449, n466, n483, n500, n501, n518, n535,
    n552;
  assign n265 = ~count[4]  & ~count[5] ;
  assign n266 = ~count[6]  & count[7] ;
  assign n267 = n265 & n266;
  assign n268 = ~count[0]  & ~count[2] ;
  assign n269 = ~count[1]  & ~count[3] ;
  assign n270 = n268 & n269;
  assign selectp1[0]  = n267 & n270;
  assign n272 = count[0]  & ~count[2] ;
  assign n273 = n269 & n272;
  assign selectp1[1]  = n267 & n273;
  assign n275 = count[1]  & ~count[3] ;
  assign n276 = n268 & n275;
  assign selectp1[2]  = n267 & n276;
  assign n278 = n272 & n275;
  assign selectp1[3]  = n267 & n278;
  assign n280 = ~count[0]  & count[2] ;
  assign n281 = n269 & n280;
  assign selectp1[4]  = n267 & n281;
  assign n283 = count[0]  & count[2] ;
  assign n284 = n269 & n283;
  assign selectp1[5]  = n267 & n284;
  assign n286 = n275 & n280;
  assign selectp1[6]  = n267 & n286;
  assign n288 = n275 & n283;
  assign selectp1[7]  = n267 & n288;
  assign n290 = ~count[1]  & count[3] ;
  assign n291 = n268 & n290;
  assign selectp1[8]  = n267 & n291;
  assign n293 = n272 & n290;
  assign selectp1[9]  = n267 & n293;
  assign n295 = count[1]  & count[3] ;
  assign n296 = n268 & n295;
  assign selectp1[10]  = n267 & n296;
  assign n298 = n272 & n295;
  assign selectp1[11]  = n267 & n298;
  assign n300 = n280 & n290;
  assign selectp1[12]  = n267 & n300;
  assign n302 = n283 & n290;
  assign selectp1[13]  = n267 & n302;
  assign n304 = n280 & n295;
  assign selectp1[14]  = n267 & n304;
  assign n306 = n283 & n295;
  assign selectp1[15]  = n267 & n306;
  assign n308 = count[4]  & ~count[5] ;
  assign n309 = n266 & n308;
  assign selectp1[16]  = n270 & n309;
  assign selectp1[17]  = n273 & n309;
  assign selectp1[18]  = n276 & n309;
  assign selectp1[19]  = n278 & n309;
  assign selectp1[20]  = n281 & n309;
  assign selectp1[21]  = n284 & n309;
  assign selectp1[22]  = n286 & n309;
  assign selectp1[23]  = n288 & n309;
  assign selectp1[24]  = n291 & n309;
  assign selectp1[25]  = n293 & n309;
  assign selectp1[26]  = n296 & n309;
  assign selectp1[27]  = n298 & n309;
  assign selectp1[28]  = n300 & n309;
  assign selectp1[29]  = n302 & n309;
  assign selectp1[30]  = n304 & n309;
  assign selectp1[31]  = n306 & n309;
  assign n326 = ~count[4]  & count[5] ;
  assign n327 = n266 & n326;
  assign selectp1[32]  = n270 & n327;
  assign selectp1[33]  = n273 & n327;
  assign selectp1[34]  = n276 & n327;
  assign selectp1[35]  = n278 & n327;
  assign selectp1[36]  = n281 & n327;
  assign selectp1[37]  = n284 & n327;
  assign selectp1[38]  = n286 & n327;
  assign selectp1[39]  = n288 & n327;
  assign selectp1[40]  = n291 & n327;
  assign selectp1[41]  = n293 & n327;
  assign selectp1[42]  = n296 & n327;
  assign selectp1[43]  = n298 & n327;
  assign selectp1[44]  = n300 & n327;
  assign selectp1[45]  = n302 & n327;
  assign selectp1[46]  = n304 & n327;
  assign selectp1[47]  = n306 & n327;
  assign n344 = count[4]  & count[5] ;
  assign n345 = n266 & n344;
  assign selectp1[48]  = n270 & n345;
  assign selectp1[49]  = n273 & n345;
  assign selectp1[50]  = n276 & n345;
  assign selectp1[51]  = n278 & n345;
  assign selectp1[52]  = n281 & n345;
  assign selectp1[53]  = n284 & n345;
  assign selectp1[54]  = n286 & n345;
  assign selectp1[55]  = n288 & n345;
  assign selectp1[56]  = n291 & n345;
  assign selectp1[57]  = n293 & n345;
  assign selectp1[58]  = n296 & n345;
  assign selectp1[59]  = n298 & n345;
  assign selectp1[60]  = n300 & n345;
  assign selectp1[61]  = n302 & n345;
  assign selectp1[62]  = n304 & n345;
  assign selectp1[63]  = n306 & n345;
  assign n362 = count[6]  & count[7] ;
  assign n363 = n265 & n362;
  assign selectp1[64]  = n270 & n363;
  assign selectp1[65]  = n273 & n363;
  assign selectp1[66]  = n276 & n363;
  assign selectp1[67]  = n278 & n363;
  assign selectp1[68]  = n281 & n363;
  assign selectp1[69]  = n284 & n363;
  assign selectp1[70]  = n286 & n363;
  assign selectp1[71]  = n288 & n363;
  assign selectp1[72]  = n291 & n363;
  assign selectp1[73]  = n293 & n363;
  assign selectp1[74]  = n296 & n363;
  assign selectp1[75]  = n298 & n363;
  assign selectp1[76]  = n300 & n363;
  assign selectp1[77]  = n302 & n363;
  assign selectp1[78]  = n304 & n363;
  assign selectp1[79]  = n306 & n363;
  assign n380 = n308 & n362;
  assign selectp1[80]  = n270 & n380;
  assign selectp1[81]  = n273 & n380;
  assign selectp1[82]  = n276 & n380;
  assign selectp1[83]  = n278 & n380;
  assign selectp1[84]  = n281 & n380;
  assign selectp1[85]  = n284 & n380;
  assign selectp1[86]  = n286 & n380;
  assign selectp1[87]  = n288 & n380;
  assign selectp1[88]  = n291 & n380;
  assign selectp1[89]  = n293 & n380;
  assign selectp1[90]  = n296 & n380;
  assign selectp1[91]  = n298 & n380;
  assign selectp1[92]  = n300 & n380;
  assign selectp1[93]  = n302 & n380;
  assign selectp1[94]  = n304 & n380;
  assign selectp1[95]  = n306 & n380;
  assign n397 = n326 & n362;
  assign selectp1[96]  = n270 & n397;
  assign selectp1[97]  = n273 & n397;
  assign selectp1[98]  = n276 & n397;
  assign selectp1[99]  = n278 & n397;
  assign selectp1[100]  = n281 & n397;
  assign selectp1[101]  = n284 & n397;
  assign selectp1[102]  = n286 & n397;
  assign selectp1[103]  = n288 & n397;
  assign selectp1[104]  = n291 & n397;
  assign selectp1[105]  = n293 & n397;
  assign selectp1[106]  = n296 & n397;
  assign selectp1[107]  = n298 & n397;
  assign selectp1[108]  = n300 & n397;
  assign selectp1[109]  = n302 & n397;
  assign selectp1[110]  = n304 & n397;
  assign selectp1[111]  = n306 & n397;
  assign n414 = n344 & n362;
  assign selectp1[112]  = n270 & n414;
  assign selectp1[113]  = n273 & n414;
  assign selectp1[114]  = n276 & n414;
  assign selectp1[115]  = n278 & n414;
  assign selectp1[116]  = n281 & n414;
  assign selectp1[117]  = n284 & n414;
  assign selectp1[118]  = n286 & n414;
  assign selectp1[119]  = n288 & n414;
  assign selectp1[120]  = n291 & n414;
  assign selectp1[121]  = n293 & n414;
  assign selectp1[122]  = n296 & n414;
  assign selectp1[123]  = n298 & n414;
  assign selectp1[124]  = n300 & n414;
  assign selectp1[125]  = n302 & n414;
  assign selectp1[126]  = n304 & n414;
  assign selectp1[127]  = n306 & n414;
  assign n431 = ~count[6]  & ~count[7] ;
  assign n432 = n265 & n431;
  assign selectp2[0]  = n270 & n432;
  assign selectp2[1]  = n273 & n432;
  assign selectp2[2]  = n276 & n432;
  assign selectp2[3]  = n278 & n432;
  assign selectp2[4]  = n281 & n432;
  assign selectp2[5]  = n284 & n432;
  assign selectp2[6]  = n286 & n432;
  assign selectp2[7]  = n288 & n432;
  assign selectp2[8]  = n291 & n432;
  assign selectp2[9]  = n293 & n432;
  assign selectp2[10]  = n296 & n432;
  assign selectp2[11]  = n298 & n432;
  assign selectp2[12]  = n300 & n432;
  assign selectp2[13]  = n302 & n432;
  assign selectp2[14]  = n304 & n432;
  assign selectp2[15]  = n306 & n432;
  assign n449 = n308 & n431;
  assign selectp2[16]  = n270 & n449;
  assign selectp2[17]  = n273 & n449;
  assign selectp2[18]  = n276 & n449;
  assign selectp2[19]  = n278 & n449;
  assign selectp2[20]  = n281 & n449;
  assign selectp2[21]  = n284 & n449;
  assign selectp2[22]  = n286 & n449;
  assign selectp2[23]  = n288 & n449;
  assign selectp2[24]  = n291 & n449;
  assign selectp2[25]  = n293 & n449;
  assign selectp2[26]  = n296 & n449;
  assign selectp2[27]  = n298 & n449;
  assign selectp2[28]  = n300 & n449;
  assign selectp2[29]  = n302 & n449;
  assign selectp2[30]  = n304 & n449;
  assign selectp2[31]  = n306 & n449;
  assign n466 = n326 & n431;
  assign selectp2[32]  = n270 & n466;
  assign selectp2[33]  = n273 & n466;
  assign selectp2[34]  = n276 & n466;
  assign selectp2[35]  = n278 & n466;
  assign selectp2[36]  = n281 & n466;
  assign selectp2[37]  = n284 & n466;
  assign selectp2[38]  = n286 & n466;
  assign selectp2[39]  = n288 & n466;
  assign selectp2[40]  = n291 & n466;
  assign selectp2[41]  = n293 & n466;
  assign selectp2[42]  = n296 & n466;
  assign selectp2[43]  = n298 & n466;
  assign selectp2[44]  = n300 & n466;
  assign selectp2[45]  = n302 & n466;
  assign selectp2[46]  = n304 & n466;
  assign selectp2[47]  = n306 & n466;
  assign n483 = n344 & n431;
  assign selectp2[48]  = n270 & n483;
  assign selectp2[49]  = n273 & n483;
  assign selectp2[50]  = n276 & n483;
  assign selectp2[51]  = n278 & n483;
  assign selectp2[52]  = n281 & n483;
  assign selectp2[53]  = n284 & n483;
  assign selectp2[54]  = n286 & n483;
  assign selectp2[55]  = n288 & n483;
  assign selectp2[56]  = n291 & n483;
  assign selectp2[57]  = n293 & n483;
  assign selectp2[58]  = n296 & n483;
  assign selectp2[59]  = n298 & n483;
  assign selectp2[60]  = n300 & n483;
  assign selectp2[61]  = n302 & n483;
  assign selectp2[62]  = n304 & n483;
  assign selectp2[63]  = n306 & n483;
  assign n500 = count[6]  & ~count[7] ;
  assign n501 = n265 & n500;
  assign selectp2[64]  = n270 & n501;
  assign selectp2[65]  = n273 & n501;
  assign selectp2[66]  = n276 & n501;
  assign selectp2[67]  = n278 & n501;
  assign selectp2[68]  = n281 & n501;
  assign selectp2[69]  = n284 & n501;
  assign selectp2[70]  = n286 & n501;
  assign selectp2[71]  = n288 & n501;
  assign selectp2[72]  = n291 & n501;
  assign selectp2[73]  = n293 & n501;
  assign selectp2[74]  = n296 & n501;
  assign selectp2[75]  = n298 & n501;
  assign selectp2[76]  = n300 & n501;
  assign selectp2[77]  = n302 & n501;
  assign selectp2[78]  = n304 & n501;
  assign selectp2[79]  = n306 & n501;
  assign n518 = n308 & n500;
  assign selectp2[80]  = n270 & n518;
  assign selectp2[81]  = n273 & n518;
  assign selectp2[82]  = n276 & n518;
  assign selectp2[83]  = n278 & n518;
  assign selectp2[84]  = n281 & n518;
  assign selectp2[85]  = n284 & n518;
  assign selectp2[86]  = n286 & n518;
  assign selectp2[87]  = n288 & n518;
  assign selectp2[88]  = n291 & n518;
  assign selectp2[89]  = n293 & n518;
  assign selectp2[90]  = n296 & n518;
  assign selectp2[91]  = n298 & n518;
  assign selectp2[92]  = n300 & n518;
  assign selectp2[93]  = n302 & n518;
  assign selectp2[94]  = n304 & n518;
  assign selectp2[95]  = n306 & n518;
  assign n535 = n326 & n500;
  assign selectp2[96]  = n270 & n535;
  assign selectp2[97]  = n273 & n535;
  assign selectp2[98]  = n276 & n535;
  assign selectp2[99]  = n278 & n535;
  assign selectp2[100]  = n281 & n535;
  assign selectp2[101]  = n284 & n535;
  assign selectp2[102]  = n286 & n535;
  assign selectp2[103]  = n288 & n535;
  assign selectp2[104]  = n291 & n535;
  assign selectp2[105]  = n293 & n535;
  assign selectp2[106]  = n296 & n535;
  assign selectp2[107]  = n298 & n535;
  assign selectp2[108]  = n300 & n535;
  assign selectp2[109]  = n302 & n535;
  assign selectp2[110]  = n304 & n535;
  assign selectp2[111]  = n306 & n535;
  assign n552 = n344 & n500;
  assign selectp2[112]  = n270 & n552;
  assign selectp2[113]  = n273 & n552;
  assign selectp2[114]  = n276 & n552;
  assign selectp2[115]  = n278 & n552;
  assign selectp2[116]  = n281 & n552;
  assign selectp2[117]  = n284 & n552;
  assign selectp2[118]  = n286 & n552;
  assign selectp2[119]  = n288 & n552;
  assign selectp2[120]  = n291 & n552;
  assign selectp2[121]  = n293 & n552;
  assign selectp2[122]  = n296 & n552;
  assign selectp2[123]  = n298 & n552;
  assign selectp2[124]  = n300 & n552;
  assign selectp2[125]  = n302 & n552;
  assign selectp2[126]  = n304 & n552;
  assign selectp2[127]  = n306 & n552;
endmodule


