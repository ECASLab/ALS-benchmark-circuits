

`timescale 1ns/1ps


//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:28:18 08/24/2011 
// Design Name: 
// Module Name:    q15_add 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module qadd #(parameter Q = 15, N = 32)
	(
    input [N-1:0] a,
    input [N-1:0] b,
    output [N-1:0] c
    );

reg [N-1:0] res;

assign c = res;

always @(a,b) begin
	// both negative or both positive
	if(a[N-1] == b[N-1]) begin						//	Since they have the same sign, absolute magnitude increases
		res[N-2:0] = a[N-2:0] + b[N-2:0];		//		So we just add the two numbers
		res[N-1] = a[N-1];							//		and set the sign appropriately...  Doesn't matter which one we use, 
															//		they both have the same sign
															//	Do the sign last, on the off-chance there was an overflow...  
		end												//		Not doing any error checking on this...
	//	one of them is negative...
	else if(a[N-1] == 0 && b[N-1] == 1) begin		//	subtract a-b
		if( a[N-2:0] > b[N-2:0] ) begin					//	if a is greater than b,
			res[N-2:0] = a[N-2:0] - b[N-2:0];			//		then just subtract b from a
			res[N-1] = 0;										//		and manually set the sign to positive
			end
		else begin												//	if a is less than b,
			res[N-2:0] = b[N-2:0] - a[N-2:0];			//		we'll actually subtract a from b to avoid a 2's complement answer
			if (res[N-2:0] == 0)
				res[N-1] = 0;										//		I don't like negative zero....
			else
				res[N-1] = 1;										//		and manually set the sign to negative
			end
		end
	else begin												//	subtract b-a (a negative, b positive)
		if( a[N-2:0] > b[N-2:0] ) begin					//	if a is greater than b,
			res[N-2:0] = a[N-2:0] - b[N-2:0];			//		we'll actually subtract b from a to avoid a 2's complement answer
			if (res[N-2:0] == 0)
				res[N-1] = 0;										//		I don't like negative zero....
			else
				res[N-1] = 1;										//		and manually set the sign to negative
			end
		else begin												//	if a is less than b,
			res[N-2:0] = b[N-2:0] - a[N-2:0];			//		then just subtract a from b
			res[N-1] = 0;										//		and manually set the sign to positive
			end
		end
	end
endmodule

module qmult #(parameter Q=15, N=32)
	(i_multiplicand,i_multiplier,o_result,ovr);
	 input	[N-1:0]	i_multiplicand;
	 input	[N-1:0]	i_multiplier;
	 output	[N-1:0]	o_result;
	 //	The underlying assumption, here, is that both fixed-point values are of the same length (N,Q)
	 //		Because of this, the results will be of length N+N = 2N bits....
	 //		This also simplifies the hand-back of results, as the binimal point 
	 //		will always be in the same location...
	output reg ovr;
	wire [2*N-1:0] r_result;		//	Multiplication by 2 values of N bits requires a register that is N+N = 2N deep...
	wire [N-1:0] r_RetVal;
	
//--------------------------------------------------------------------------------
	assign o_result = r_RetVal;	//Only handing back the same number of bits as we received...with fixed point in same location...
	assign r_RetVal[N-1] = i_multiplicand[N-1] ^ i_multiplier[N-1];
	assign r_RetVal[N-2:0] = r_result[N-2+Q:Q];
//---------------------------------------------------------------------------------

        always @(r_result) begin	
		if (r_result[2*N-2:N-1+Q] > 0)	
			ovr = 1'b1;
		else
			ovr = 1'b0;
		
	end

	Multiplier_31_0_3000 mul0 (r_result, {1'b0,i_multiplicand[N-2:0]}, {1'b0,i_multiplier[N-2:0]});
	

endmodule

/*----------------------------------------------------------------------------
  Copyright (c) 2004 Aoki laboratory. All rights reserved.

  Top module: Multiplier_31_0_3000

  Number system: 2's complement
  Multiplicand length: 32
  Multiplier length: 32
  Partial product generation: Simple PPG
  Partial product accumulation: Wallace tree
  Final stage addition: Kogge-Stone adder
----------------------------------------------------------------------------*/

module TCDECON_31_0(TOP, R, I);
  output [30:0] R;
  output [31:31] TOP;
  input [31:0] I;
  assign TOP[31] = I[31];
  assign R[0] = I[0];
  assign R[1] = I[1];
  assign R[2] = I[2];
  assign R[3] = I[3];
  assign R[4] = I[4];
  assign R[5] = I[5];
  assign R[6] = I[6];
  assign R[7] = I[7];
  assign R[8] = I[8];
  assign R[9] = I[9];
  assign R[10] = I[10];
  assign R[11] = I[11];
  assign R[12] = I[12];
  assign R[13] = I[13];
  assign R[14] = I[14];
  assign R[15] = I[15];
  assign R[16] = I[16];
  assign R[17] = I[17];
  assign R[18] = I[18];
  assign R[19] = I[19];
  assign R[20] = I[20];
  assign R[21] = I[21];
  assign R[22] = I[22];
  assign R[23] = I[23];
  assign R[24] = I[24];
  assign R[25] = I[25];
  assign R[26] = I[26];
  assign R[27] = I[27];
  assign R[28] = I[28];
  assign R[29] = I[29];
  assign R[30] = I[30];
endmodule

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule


module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_31(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_32(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_33(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_34(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_35(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_36(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_37(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_38(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_39(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_40(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_41(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_42(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_43(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_44(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_45(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_46(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_47(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_48(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_49(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_50(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_51(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_52(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_53(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_54(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_55(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_56(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_57(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_58(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_59(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_60(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_61(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UN1BPPG_0_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_1_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_2_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_3_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_4_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_5_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_6_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_7_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_8_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_9_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_10_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_11_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_12_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_13_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_14_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_15_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_16_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_17_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_18_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_19_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_20_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_21_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_22_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_23_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_24_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_25_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_26_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_27_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_28_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_29_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_30_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUB1BPPG_31_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBOne_32(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_32(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_28(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_29(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_30(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_31(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_32(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_33(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_33(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_34(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_35(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_36(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_35(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_36(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_37(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_38(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_39(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_38(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_39(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_40(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_41(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_42(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_34(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_35(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_37(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_39(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_41(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_42(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_43(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_14(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_43(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_44(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_45(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_46(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_17(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_45(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_46(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_47(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_48(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_49(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_20(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_48(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_49(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_50(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_51(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_52(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_23(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_51(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_52(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_53(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_54(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_55(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_26(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_54(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_55(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_56(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_57(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_58(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_29(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_57(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_58(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_59(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_60(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_61(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_36(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_37(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_38(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_42(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_43(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_15(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_47(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_48(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_19(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_50(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_52(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_24(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_56(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_57(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_28(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_59(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_61(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_40(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_41(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_13(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_46(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_47(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_21(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_53(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_54(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_27(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_58(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_62(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_44(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_45(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_18(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_49(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_30(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_60(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_61(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_62(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_50(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_51(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_53(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_25(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_56(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_62(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_63(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_16(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_55(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_59(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_60(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_22(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_63(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBZero_64_64(O);
  output [64:64] O;
  assign O[64] = 0;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriKSA_64_9(S, X, Y, Cin);
  output [65:9] S;
  input Cin;
  input [64:9] X;
  input [64:9] Y;
  wire [64:9] G0;
  wire [64:9] G1;
  wire [64:9] G2;
  wire [64:9] G3;
  wire [64:9] G4;
  wire [64:9] G5;
  wire [64:9] G6;
  wire [64:9] P0;
  wire [64:9] P1;
  wire [64:9] P2;
  wire [64:9] P3;
  wire [64:9] P4;
  wire [64:9] P5;
  wire [64:9] P6;
  assign P1[9] = P0[9];
  assign G1[9] = G0[9];
  assign P2[9] = P1[9];
  assign G2[9] = G1[9];
  assign P2[10] = P1[10];
  assign G2[10] = G1[10];
  assign P3[9] = P2[9];
  assign G3[9] = G2[9];
  assign P3[10] = P2[10];
  assign G3[10] = G2[10];
  assign P3[11] = P2[11];
  assign G3[11] = G2[11];
  assign P3[12] = P2[12];
  assign G3[12] = G2[12];
  assign P4[9] = P3[9];
  assign G4[9] = G3[9];
  assign P4[10] = P3[10];
  assign G4[10] = G3[10];
  assign P4[11] = P3[11];
  assign G4[11] = G3[11];
  assign P4[12] = P3[12];
  assign G4[12] = G3[12];
  assign P4[13] = P3[13];
  assign G4[13] = G3[13];
  assign P4[14] = P3[14];
  assign G4[14] = G3[14];
  assign P4[15] = P3[15];
  assign G4[15] = G3[15];
  assign P4[16] = P3[16];
  assign G4[16] = G3[16];
  assign P5[9] = P4[9];
  assign G5[9] = G4[9];
  assign P5[10] = P4[10];
  assign G5[10] = G4[10];
  assign P5[11] = P4[11];
  assign G5[11] = G4[11];
  assign P5[12] = P4[12];
  assign G5[12] = G4[12];
  assign P5[13] = P4[13];
  assign G5[13] = G4[13];
  assign P5[14] = P4[14];
  assign G5[14] = G4[14];
  assign P5[15] = P4[15];
  assign G5[15] = G4[15];
  assign P5[16] = P4[16];
  assign G5[16] = G4[16];
  assign P5[17] = P4[17];
  assign G5[17] = G4[17];
  assign P5[18] = P4[18];
  assign G5[18] = G4[18];
  assign P5[19] = P4[19];
  assign G5[19] = G4[19];
  assign P5[20] = P4[20];
  assign G5[20] = G4[20];
  assign P5[21] = P4[21];
  assign G5[21] = G4[21];
  assign P5[22] = P4[22];
  assign G5[22] = G4[22];
  assign P5[23] = P4[23];
  assign G5[23] = G4[23];
  assign P5[24] = P4[24];
  assign G5[24] = G4[24];
  assign P6[9] = P5[9];
  assign G6[9] = G5[9];
  assign P6[10] = P5[10];
  assign G6[10] = G5[10];
  assign P6[11] = P5[11];
  assign G6[11] = G5[11];
  assign P6[12] = P5[12];
  assign G6[12] = G5[12];
  assign P6[13] = P5[13];
  assign G6[13] = G5[13];
  assign P6[14] = P5[14];
  assign G6[14] = G5[14];
  assign P6[15] = P5[15];
  assign G6[15] = G5[15];
  assign P6[16] = P5[16];
  assign G6[16] = G5[16];
  assign P6[17] = P5[17];
  assign G6[17] = G5[17];
  assign P6[18] = P5[18];
  assign G6[18] = G5[18];
  assign P6[19] = P5[19];
  assign G6[19] = G5[19];
  assign P6[20] = P5[20];
  assign G6[20] = G5[20];
  assign P6[21] = P5[21];
  assign G6[21] = G5[21];
  assign P6[22] = P5[22];
  assign G6[22] = G5[22];
  assign P6[23] = P5[23];
  assign G6[23] = G5[23];
  assign P6[24] = P5[24];
  assign G6[24] = G5[24];
  assign P6[25] = P5[25];
  assign G6[25] = G5[25];
  assign P6[26] = P5[26];
  assign G6[26] = G5[26];
  assign P6[27] = P5[27];
  assign G6[27] = G5[27];
  assign P6[28] = P5[28];
  assign G6[28] = G5[28];
  assign P6[29] = P5[29];
  assign G6[29] = G5[29];
  assign P6[30] = P5[30];
  assign G6[30] = G5[30];
  assign P6[31] = P5[31];
  assign G6[31] = G5[31];
  assign P6[32] = P5[32];
  assign G6[32] = G5[32];
  assign P6[33] = P5[33];
  assign G6[33] = G5[33];
  assign P6[34] = P5[34];
  assign G6[34] = G5[34];
  assign P6[35] = P5[35];
  assign G6[35] = G5[35];
  assign P6[36] = P5[36];
  assign G6[36] = G5[36];
  assign P6[37] = P5[37];
  assign G6[37] = G5[37];
  assign P6[38] = P5[38];
  assign G6[38] = G5[38];
  assign P6[39] = P5[39];
  assign G6[39] = G5[39];
  assign P6[40] = P5[40];
  assign G6[40] = G5[40];
  assign S[9] = Cin ^ P0[9];
  assign S[10] = ( G6[9] | ( P6[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G6[10] | ( P6[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G6[11] | ( P6[11] & Cin ) ) ^ P0[12];
  assign S[13] = ( G6[12] | ( P6[12] & Cin ) ) ^ P0[13];
  assign S[14] = ( G6[13] | ( P6[13] & Cin ) ) ^ P0[14];
  assign S[15] = ( G6[14] | ( P6[14] & Cin ) ) ^ P0[15];
  assign S[16] = ( G6[15] | ( P6[15] & Cin ) ) ^ P0[16];
  assign S[17] = ( G6[16] | ( P6[16] & Cin ) ) ^ P0[17];
  assign S[18] = ( G6[17] | ( P6[17] & Cin ) ) ^ P0[18];
  assign S[19] = ( G6[18] | ( P6[18] & Cin ) ) ^ P0[19];
  assign S[20] = ( G6[19] | ( P6[19] & Cin ) ) ^ P0[20];
  assign S[21] = ( G6[20] | ( P6[20] & Cin ) ) ^ P0[21];
  assign S[22] = ( G6[21] | ( P6[21] & Cin ) ) ^ P0[22];
  assign S[23] = ( G6[22] | ( P6[22] & Cin ) ) ^ P0[23];
  assign S[24] = ( G6[23] | ( P6[23] & Cin ) ) ^ P0[24];
  assign S[25] = ( G6[24] | ( P6[24] & Cin ) ) ^ P0[25];
  assign S[26] = ( G6[25] | ( P6[25] & Cin ) ) ^ P0[26];
  assign S[27] = ( G6[26] | ( P6[26] & Cin ) ) ^ P0[27];
  assign S[28] = ( G6[27] | ( P6[27] & Cin ) ) ^ P0[28];
  assign S[29] = ( G6[28] | ( P6[28] & Cin ) ) ^ P0[29];
  assign S[30] = ( G6[29] | ( P6[29] & Cin ) ) ^ P0[30];
  assign S[31] = ( G6[30] | ( P6[30] & Cin ) ) ^ P0[31];
  assign S[32] = ( G6[31] | ( P6[31] & Cin ) ) ^ P0[32];
  assign S[33] = ( G6[32] | ( P6[32] & Cin ) ) ^ P0[33];
  assign S[34] = ( G6[33] | ( P6[33] & Cin ) ) ^ P0[34];
  assign S[35] = ( G6[34] | ( P6[34] & Cin ) ) ^ P0[35];
  assign S[36] = ( G6[35] | ( P6[35] & Cin ) ) ^ P0[36];
  assign S[37] = ( G6[36] | ( P6[36] & Cin ) ) ^ P0[37];
  assign S[38] = ( G6[37] | ( P6[37] & Cin ) ) ^ P0[38];
  assign S[39] = ( G6[38] | ( P6[38] & Cin ) ) ^ P0[39];
  assign S[40] = ( G6[39] | ( P6[39] & Cin ) ) ^ P0[40];
  assign S[41] = ( G6[40] | ( P6[40] & Cin ) ) ^ P0[41];
  assign S[42] = ( G6[41] | ( P6[41] & Cin ) ) ^ P0[42];
  assign S[43] = ( G6[42] | ( P6[42] & Cin ) ) ^ P0[43];
  assign S[44] = ( G6[43] | ( P6[43] & Cin ) ) ^ P0[44];
  assign S[45] = ( G6[44] | ( P6[44] & Cin ) ) ^ P0[45];
  assign S[46] = ( G6[45] | ( P6[45] & Cin ) ) ^ P0[46];
  assign S[47] = ( G6[46] | ( P6[46] & Cin ) ) ^ P0[47];
  assign S[48] = ( G6[47] | ( P6[47] & Cin ) ) ^ P0[48];
  assign S[49] = ( G6[48] | ( P6[48] & Cin ) ) ^ P0[49];
  assign S[50] = ( G6[49] | ( P6[49] & Cin ) ) ^ P0[50];
  assign S[51] = ( G6[50] | ( P6[50] & Cin ) ) ^ P0[51];
  assign S[52] = ( G6[51] | ( P6[51] & Cin ) ) ^ P0[52];
  assign S[53] = ( G6[52] | ( P6[52] & Cin ) ) ^ P0[53];
  assign S[54] = ( G6[53] | ( P6[53] & Cin ) ) ^ P0[54];
  assign S[55] = ( G6[54] | ( P6[54] & Cin ) ) ^ P0[55];
  assign S[56] = ( G6[55] | ( P6[55] & Cin ) ) ^ P0[56];
  assign S[57] = ( G6[56] | ( P6[56] & Cin ) ) ^ P0[57];
  assign S[58] = ( G6[57] | ( P6[57] & Cin ) ) ^ P0[58];
  assign S[59] = ( G6[58] | ( P6[58] & Cin ) ) ^ P0[59];
  assign S[60] = ( G6[59] | ( P6[59] & Cin ) ) ^ P0[60];
  assign S[61] = ( G6[60] | ( P6[60] & Cin ) ) ^ P0[61];
  assign S[62] = ( G6[61] | ( P6[61] & Cin ) ) ^ P0[62];
  assign S[63] = ( G6[62] | ( P6[62] & Cin ) ) ^ P0[63];
  assign S[64] = ( G6[63] | ( P6[63] & Cin ) ) ^ P0[64];
  assign S[65] = G6[64] | ( P6[64] & Cin );
  GPGenerator U0 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U1 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U2 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U3 (G0[12], P0[12], X[12], Y[12]);
  GPGenerator U4 (G0[13], P0[13], X[13], Y[13]);
  GPGenerator U5 (G0[14], P0[14], X[14], Y[14]);
  GPGenerator U6 (G0[15], P0[15], X[15], Y[15]);
  GPGenerator U7 (G0[16], P0[16], X[16], Y[16]);
  GPGenerator U8 (G0[17], P0[17], X[17], Y[17]);
  GPGenerator U9 (G0[18], P0[18], X[18], Y[18]);
  GPGenerator U10 (G0[19], P0[19], X[19], Y[19]);
  GPGenerator U11 (G0[20], P0[20], X[20], Y[20]);
  GPGenerator U12 (G0[21], P0[21], X[21], Y[21]);
  GPGenerator U13 (G0[22], P0[22], X[22], Y[22]);
  GPGenerator U14 (G0[23], P0[23], X[23], Y[23]);
  GPGenerator U15 (G0[24], P0[24], X[24], Y[24]);
  GPGenerator U16 (G0[25], P0[25], X[25], Y[25]);
  GPGenerator U17 (G0[26], P0[26], X[26], Y[26]);
  GPGenerator U18 (G0[27], P0[27], X[27], Y[27]);
  GPGenerator U19 (G0[28], P0[28], X[28], Y[28]);
  GPGenerator U20 (G0[29], P0[29], X[29], Y[29]);
  GPGenerator U21 (G0[30], P0[30], X[30], Y[30]);
  GPGenerator U22 (G0[31], P0[31], X[31], Y[31]);
  GPGenerator U23 (G0[32], P0[32], X[32], Y[32]);
  GPGenerator U24 (G0[33], P0[33], X[33], Y[33]);
  GPGenerator U25 (G0[34], P0[34], X[34], Y[34]);
  GPGenerator U26 (G0[35], P0[35], X[35], Y[35]);
  GPGenerator U27 (G0[36], P0[36], X[36], Y[36]);
  GPGenerator U28 (G0[37], P0[37], X[37], Y[37]);
  GPGenerator U29 (G0[38], P0[38], X[38], Y[38]);
  GPGenerator U30 (G0[39], P0[39], X[39], Y[39]);
  GPGenerator U31 (G0[40], P0[40], X[40], Y[40]);
  GPGenerator U32 (G0[41], P0[41], X[41], Y[41]);
  GPGenerator U33 (G0[42], P0[42], X[42], Y[42]);
  GPGenerator U34 (G0[43], P0[43], X[43], Y[43]);
  GPGenerator U35 (G0[44], P0[44], X[44], Y[44]);
  GPGenerator U36 (G0[45], P0[45], X[45], Y[45]);
  GPGenerator U37 (G0[46], P0[46], X[46], Y[46]);
  GPGenerator U38 (G0[47], P0[47], X[47], Y[47]);
  GPGenerator U39 (G0[48], P0[48], X[48], Y[48]);
  GPGenerator U40 (G0[49], P0[49], X[49], Y[49]);
  GPGenerator U41 (G0[50], P0[50], X[50], Y[50]);
  GPGenerator U42 (G0[51], P0[51], X[51], Y[51]);
  GPGenerator U43 (G0[52], P0[52], X[52], Y[52]);
  GPGenerator U44 (G0[53], P0[53], X[53], Y[53]);
  GPGenerator U45 (G0[54], P0[54], X[54], Y[54]);
  GPGenerator U46 (G0[55], P0[55], X[55], Y[55]);
  GPGenerator U47 (G0[56], P0[56], X[56], Y[56]);
  GPGenerator U48 (G0[57], P0[57], X[57], Y[57]);
  GPGenerator U49 (G0[58], P0[58], X[58], Y[58]);
  GPGenerator U50 (G0[59], P0[59], X[59], Y[59]);
  GPGenerator U51 (G0[60], P0[60], X[60], Y[60]);
  GPGenerator U52 (G0[61], P0[61], X[61], Y[61]);
  GPGenerator U53 (G0[62], P0[62], X[62], Y[62]);
  GPGenerator U54 (G0[63], P0[63], X[63], Y[63]);
  GPGenerator U55 (G0[64], P0[64], X[64], Y[64]);
  CarryOperator U56 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U57 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U58 (G1[12], P1[12], G0[12], P0[12], G0[11], P0[11]);
  CarryOperator U59 (G1[13], P1[13], G0[13], P0[13], G0[12], P0[12]);
  CarryOperator U60 (G1[14], P1[14], G0[14], P0[14], G0[13], P0[13]);
  CarryOperator U61 (G1[15], P1[15], G0[15], P0[15], G0[14], P0[14]);
  CarryOperator U62 (G1[16], P1[16], G0[16], P0[16], G0[15], P0[15]);
  CarryOperator U63 (G1[17], P1[17], G0[17], P0[17], G0[16], P0[16]);
  CarryOperator U64 (G1[18], P1[18], G0[18], P0[18], G0[17], P0[17]);
  CarryOperator U65 (G1[19], P1[19], G0[19], P0[19], G0[18], P0[18]);
  CarryOperator U66 (G1[20], P1[20], G0[20], P0[20], G0[19], P0[19]);
  CarryOperator U67 (G1[21], P1[21], G0[21], P0[21], G0[20], P0[20]);
  CarryOperator U68 (G1[22], P1[22], G0[22], P0[22], G0[21], P0[21]);
  CarryOperator U69 (G1[23], P1[23], G0[23], P0[23], G0[22], P0[22]);
  CarryOperator U70 (G1[24], P1[24], G0[24], P0[24], G0[23], P0[23]);
  CarryOperator U71 (G1[25], P1[25], G0[25], P0[25], G0[24], P0[24]);
  CarryOperator U72 (G1[26], P1[26], G0[26], P0[26], G0[25], P0[25]);
  CarryOperator U73 (G1[27], P1[27], G0[27], P0[27], G0[26], P0[26]);
  CarryOperator U74 (G1[28], P1[28], G0[28], P0[28], G0[27], P0[27]);
  CarryOperator U75 (G1[29], P1[29], G0[29], P0[29], G0[28], P0[28]);
  CarryOperator U76 (G1[30], P1[30], G0[30], P0[30], G0[29], P0[29]);
  CarryOperator U77 (G1[31], P1[31], G0[31], P0[31], G0[30], P0[30]);
  CarryOperator U78 (G1[32], P1[32], G0[32], P0[32], G0[31], P0[31]);
  CarryOperator U79 (G1[33], P1[33], G0[33], P0[33], G0[32], P0[32]);
  CarryOperator U80 (G1[34], P1[34], G0[34], P0[34], G0[33], P0[33]);
  CarryOperator U81 (G1[35], P1[35], G0[35], P0[35], G0[34], P0[34]);
  CarryOperator U82 (G1[36], P1[36], G0[36], P0[36], G0[35], P0[35]);
  CarryOperator U83 (G1[37], P1[37], G0[37], P0[37], G0[36], P0[36]);
  CarryOperator U84 (G1[38], P1[38], G0[38], P0[38], G0[37], P0[37]);
  CarryOperator U85 (G1[39], P1[39], G0[39], P0[39], G0[38], P0[38]);
  CarryOperator U86 (G1[40], P1[40], G0[40], P0[40], G0[39], P0[39]);
  CarryOperator U87 (G1[41], P1[41], G0[41], P0[41], G0[40], P0[40]);
  CarryOperator U88 (G1[42], P1[42], G0[42], P0[42], G0[41], P0[41]);
  CarryOperator U89 (G1[43], P1[43], G0[43], P0[43], G0[42], P0[42]);
  CarryOperator U90 (G1[44], P1[44], G0[44], P0[44], G0[43], P0[43]);
  CarryOperator U91 (G1[45], P1[45], G0[45], P0[45], G0[44], P0[44]);
  CarryOperator U92 (G1[46], P1[46], G0[46], P0[46], G0[45], P0[45]);
  CarryOperator U93 (G1[47], P1[47], G0[47], P0[47], G0[46], P0[46]);
  CarryOperator U94 (G1[48], P1[48], G0[48], P0[48], G0[47], P0[47]);
  CarryOperator U95 (G1[49], P1[49], G0[49], P0[49], G0[48], P0[48]);
  CarryOperator U96 (G1[50], P1[50], G0[50], P0[50], G0[49], P0[49]);
  CarryOperator U97 (G1[51], P1[51], G0[51], P0[51], G0[50], P0[50]);
  CarryOperator U98 (G1[52], P1[52], G0[52], P0[52], G0[51], P0[51]);
  CarryOperator U99 (G1[53], P1[53], G0[53], P0[53], G0[52], P0[52]);
  CarryOperator U100 (G1[54], P1[54], G0[54], P0[54], G0[53], P0[53]);
  CarryOperator U101 (G1[55], P1[55], G0[55], P0[55], G0[54], P0[54]);
  CarryOperator U102 (G1[56], P1[56], G0[56], P0[56], G0[55], P0[55]);
  CarryOperator U103 (G1[57], P1[57], G0[57], P0[57], G0[56], P0[56]);
  CarryOperator U104 (G1[58], P1[58], G0[58], P0[58], G0[57], P0[57]);
  CarryOperator U105 (G1[59], P1[59], G0[59], P0[59], G0[58], P0[58]);
  CarryOperator U106 (G1[60], P1[60], G0[60], P0[60], G0[59], P0[59]);
  CarryOperator U107 (G1[61], P1[61], G0[61], P0[61], G0[60], P0[60]);
  CarryOperator U108 (G1[62], P1[62], G0[62], P0[62], G0[61], P0[61]);
  CarryOperator U109 (G1[63], P1[63], G0[63], P0[63], G0[62], P0[62]);
  CarryOperator U110 (G1[64], P1[64], G0[64], P0[64], G0[63], P0[63]);
  CarryOperator U111 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U112 (G2[12], P2[12], G1[12], P1[12], G1[10], P1[10]);
  CarryOperator U113 (G2[13], P2[13], G1[13], P1[13], G1[11], P1[11]);
  CarryOperator U114 (G2[14], P2[14], G1[14], P1[14], G1[12], P1[12]);
  CarryOperator U115 (G2[15], P2[15], G1[15], P1[15], G1[13], P1[13]);
  CarryOperator U116 (G2[16], P2[16], G1[16], P1[16], G1[14], P1[14]);
  CarryOperator U117 (G2[17], P2[17], G1[17], P1[17], G1[15], P1[15]);
  CarryOperator U118 (G2[18], P2[18], G1[18], P1[18], G1[16], P1[16]);
  CarryOperator U119 (G2[19], P2[19], G1[19], P1[19], G1[17], P1[17]);
  CarryOperator U120 (G2[20], P2[20], G1[20], P1[20], G1[18], P1[18]);
  CarryOperator U121 (G2[21], P2[21], G1[21], P1[21], G1[19], P1[19]);
  CarryOperator U122 (G2[22], P2[22], G1[22], P1[22], G1[20], P1[20]);
  CarryOperator U123 (G2[23], P2[23], G1[23], P1[23], G1[21], P1[21]);
  CarryOperator U124 (G2[24], P2[24], G1[24], P1[24], G1[22], P1[22]);
  CarryOperator U125 (G2[25], P2[25], G1[25], P1[25], G1[23], P1[23]);
  CarryOperator U126 (G2[26], P2[26], G1[26], P1[26], G1[24], P1[24]);
  CarryOperator U127 (G2[27], P2[27], G1[27], P1[27], G1[25], P1[25]);
  CarryOperator U128 (G2[28], P2[28], G1[28], P1[28], G1[26], P1[26]);
  CarryOperator U129 (G2[29], P2[29], G1[29], P1[29], G1[27], P1[27]);
  CarryOperator U130 (G2[30], P2[30], G1[30], P1[30], G1[28], P1[28]);
  CarryOperator U131 (G2[31], P2[31], G1[31], P1[31], G1[29], P1[29]);
  CarryOperator U132 (G2[32], P2[32], G1[32], P1[32], G1[30], P1[30]);
  CarryOperator U133 (G2[33], P2[33], G1[33], P1[33], G1[31], P1[31]);
  CarryOperator U134 (G2[34], P2[34], G1[34], P1[34], G1[32], P1[32]);
  CarryOperator U135 (G2[35], P2[35], G1[35], P1[35], G1[33], P1[33]);
  CarryOperator U136 (G2[36], P2[36], G1[36], P1[36], G1[34], P1[34]);
  CarryOperator U137 (G2[37], P2[37], G1[37], P1[37], G1[35], P1[35]);
  CarryOperator U138 (G2[38], P2[38], G1[38], P1[38], G1[36], P1[36]);
  CarryOperator U139 (G2[39], P2[39], G1[39], P1[39], G1[37], P1[37]);
  CarryOperator U140 (G2[40], P2[40], G1[40], P1[40], G1[38], P1[38]);
  CarryOperator U141 (G2[41], P2[41], G1[41], P1[41], G1[39], P1[39]);
  CarryOperator U142 (G2[42], P2[42], G1[42], P1[42], G1[40], P1[40]);
  CarryOperator U143 (G2[43], P2[43], G1[43], P1[43], G1[41], P1[41]);
  CarryOperator U144 (G2[44], P2[44], G1[44], P1[44], G1[42], P1[42]);
  CarryOperator U145 (G2[45], P2[45], G1[45], P1[45], G1[43], P1[43]);
  CarryOperator U146 (G2[46], P2[46], G1[46], P1[46], G1[44], P1[44]);
  CarryOperator U147 (G2[47], P2[47], G1[47], P1[47], G1[45], P1[45]);
  CarryOperator U148 (G2[48], P2[48], G1[48], P1[48], G1[46], P1[46]);
  CarryOperator U149 (G2[49], P2[49], G1[49], P1[49], G1[47], P1[47]);
  CarryOperator U150 (G2[50], P2[50], G1[50], P1[50], G1[48], P1[48]);
  CarryOperator U151 (G2[51], P2[51], G1[51], P1[51], G1[49], P1[49]);
  CarryOperator U152 (G2[52], P2[52], G1[52], P1[52], G1[50], P1[50]);
  CarryOperator U153 (G2[53], P2[53], G1[53], P1[53], G1[51], P1[51]);
  CarryOperator U154 (G2[54], P2[54], G1[54], P1[54], G1[52], P1[52]);
  CarryOperator U155 (G2[55], P2[55], G1[55], P1[55], G1[53], P1[53]);
  CarryOperator U156 (G2[56], P2[56], G1[56], P1[56], G1[54], P1[54]);
  CarryOperator U157 (G2[57], P2[57], G1[57], P1[57], G1[55], P1[55]);
  CarryOperator U158 (G2[58], P2[58], G1[58], P1[58], G1[56], P1[56]);
  CarryOperator U159 (G2[59], P2[59], G1[59], P1[59], G1[57], P1[57]);
  CarryOperator U160 (G2[60], P2[60], G1[60], P1[60], G1[58], P1[58]);
  CarryOperator U161 (G2[61], P2[61], G1[61], P1[61], G1[59], P1[59]);
  CarryOperator U162 (G2[62], P2[62], G1[62], P1[62], G1[60], P1[60]);
  CarryOperator U163 (G2[63], P2[63], G1[63], P1[63], G1[61], P1[61]);
  CarryOperator U164 (G2[64], P2[64], G1[64], P1[64], G1[62], P1[62]);
  CarryOperator U165 (G3[13], P3[13], G2[13], P2[13], G2[9], P2[9]);
  CarryOperator U166 (G3[14], P3[14], G2[14], P2[14], G2[10], P2[10]);
  CarryOperator U167 (G3[15], P3[15], G2[15], P2[15], G2[11], P2[11]);
  CarryOperator U168 (G3[16], P3[16], G2[16], P2[16], G2[12], P2[12]);
  CarryOperator U169 (G3[17], P3[17], G2[17], P2[17], G2[13], P2[13]);
  CarryOperator U170 (G3[18], P3[18], G2[18], P2[18], G2[14], P2[14]);
  CarryOperator U171 (G3[19], P3[19], G2[19], P2[19], G2[15], P2[15]);
  CarryOperator U172 (G3[20], P3[20], G2[20], P2[20], G2[16], P2[16]);
  CarryOperator U173 (G3[21], P3[21], G2[21], P2[21], G2[17], P2[17]);
  CarryOperator U174 (G3[22], P3[22], G2[22], P2[22], G2[18], P2[18]);
  CarryOperator U175 (G3[23], P3[23], G2[23], P2[23], G2[19], P2[19]);
  CarryOperator U176 (G3[24], P3[24], G2[24], P2[24], G2[20], P2[20]);
  CarryOperator U177 (G3[25], P3[25], G2[25], P2[25], G2[21], P2[21]);
  CarryOperator U178 (G3[26], P3[26], G2[26], P2[26], G2[22], P2[22]);
  CarryOperator U179 (G3[27], P3[27], G2[27], P2[27], G2[23], P2[23]);
  CarryOperator U180 (G3[28], P3[28], G2[28], P2[28], G2[24], P2[24]);
  CarryOperator U181 (G3[29], P3[29], G2[29], P2[29], G2[25], P2[25]);
  CarryOperator U182 (G3[30], P3[30], G2[30], P2[30], G2[26], P2[26]);
  CarryOperator U183 (G3[31], P3[31], G2[31], P2[31], G2[27], P2[27]);
  CarryOperator U184 (G3[32], P3[32], G2[32], P2[32], G2[28], P2[28]);
  CarryOperator U185 (G3[33], P3[33], G2[33], P2[33], G2[29], P2[29]);
  CarryOperator U186 (G3[34], P3[34], G2[34], P2[34], G2[30], P2[30]);
  CarryOperator U187 (G3[35], P3[35], G2[35], P2[35], G2[31], P2[31]);
  CarryOperator U188 (G3[36], P3[36], G2[36], P2[36], G2[32], P2[32]);
  CarryOperator U189 (G3[37], P3[37], G2[37], P2[37], G2[33], P2[33]);
  CarryOperator U190 (G3[38], P3[38], G2[38], P2[38], G2[34], P2[34]);
  CarryOperator U191 (G3[39], P3[39], G2[39], P2[39], G2[35], P2[35]);
  CarryOperator U192 (G3[40], P3[40], G2[40], P2[40], G2[36], P2[36]);
  CarryOperator U193 (G3[41], P3[41], G2[41], P2[41], G2[37], P2[37]);
  CarryOperator U194 (G3[42], P3[42], G2[42], P2[42], G2[38], P2[38]);
  CarryOperator U195 (G3[43], P3[43], G2[43], P2[43], G2[39], P2[39]);
  CarryOperator U196 (G3[44], P3[44], G2[44], P2[44], G2[40], P2[40]);
  CarryOperator U197 (G3[45], P3[45], G2[45], P2[45], G2[41], P2[41]);
  CarryOperator U198 (G3[46], P3[46], G2[46], P2[46], G2[42], P2[42]);
  CarryOperator U199 (G3[47], P3[47], G2[47], P2[47], G2[43], P2[43]);
  CarryOperator U200 (G3[48], P3[48], G2[48], P2[48], G2[44], P2[44]);
  CarryOperator U201 (G3[49], P3[49], G2[49], P2[49], G2[45], P2[45]);
  CarryOperator U202 (G3[50], P3[50], G2[50], P2[50], G2[46], P2[46]);
  CarryOperator U203 (G3[51], P3[51], G2[51], P2[51], G2[47], P2[47]);
  CarryOperator U204 (G3[52], P3[52], G2[52], P2[52], G2[48], P2[48]);
  CarryOperator U205 (G3[53], P3[53], G2[53], P2[53], G2[49], P2[49]);
  CarryOperator U206 (G3[54], P3[54], G2[54], P2[54], G2[50], P2[50]);
  CarryOperator U207 (G3[55], P3[55], G2[55], P2[55], G2[51], P2[51]);
  CarryOperator U208 (G3[56], P3[56], G2[56], P2[56], G2[52], P2[52]);
  CarryOperator U209 (G3[57], P3[57], G2[57], P2[57], G2[53], P2[53]);
  CarryOperator U210 (G3[58], P3[58], G2[58], P2[58], G2[54], P2[54]);
  CarryOperator U211 (G3[59], P3[59], G2[59], P2[59], G2[55], P2[55]);
  CarryOperator U212 (G3[60], P3[60], G2[60], P2[60], G2[56], P2[56]);
  CarryOperator U213 (G3[61], P3[61], G2[61], P2[61], G2[57], P2[57]);
  CarryOperator U214 (G3[62], P3[62], G2[62], P2[62], G2[58], P2[58]);
  CarryOperator U215 (G3[63], P3[63], G2[63], P2[63], G2[59], P2[59]);
  CarryOperator U216 (G3[64], P3[64], G2[64], P2[64], G2[60], P2[60]);
  CarryOperator U217 (G4[17], P4[17], G3[17], P3[17], G3[9], P3[9]);
  CarryOperator U218 (G4[18], P4[18], G3[18], P3[18], G3[10], P3[10]);
  CarryOperator U219 (G4[19], P4[19], G3[19], P3[19], G3[11], P3[11]);
  CarryOperator U220 (G4[20], P4[20], G3[20], P3[20], G3[12], P3[12]);
  CarryOperator U221 (G4[21], P4[21], G3[21], P3[21], G3[13], P3[13]);
  CarryOperator U222 (G4[22], P4[22], G3[22], P3[22], G3[14], P3[14]);
  CarryOperator U223 (G4[23], P4[23], G3[23], P3[23], G3[15], P3[15]);
  CarryOperator U224 (G4[24], P4[24], G3[24], P3[24], G3[16], P3[16]);
  CarryOperator U225 (G4[25], P4[25], G3[25], P3[25], G3[17], P3[17]);
  CarryOperator U226 (G4[26], P4[26], G3[26], P3[26], G3[18], P3[18]);
  CarryOperator U227 (G4[27], P4[27], G3[27], P3[27], G3[19], P3[19]);
  CarryOperator U228 (G4[28], P4[28], G3[28], P3[28], G3[20], P3[20]);
  CarryOperator U229 (G4[29], P4[29], G3[29], P3[29], G3[21], P3[21]);
  CarryOperator U230 (G4[30], P4[30], G3[30], P3[30], G3[22], P3[22]);
  CarryOperator U231 (G4[31], P4[31], G3[31], P3[31], G3[23], P3[23]);
  CarryOperator U232 (G4[32], P4[32], G3[32], P3[32], G3[24], P3[24]);
  CarryOperator U233 (G4[33], P4[33], G3[33], P3[33], G3[25], P3[25]);
  CarryOperator U234 (G4[34], P4[34], G3[34], P3[34], G3[26], P3[26]);
  CarryOperator U235 (G4[35], P4[35], G3[35], P3[35], G3[27], P3[27]);
  CarryOperator U236 (G4[36], P4[36], G3[36], P3[36], G3[28], P3[28]);
  CarryOperator U237 (G4[37], P4[37], G3[37], P3[37], G3[29], P3[29]);
  CarryOperator U238 (G4[38], P4[38], G3[38], P3[38], G3[30], P3[30]);
  CarryOperator U239 (G4[39], P4[39], G3[39], P3[39], G3[31], P3[31]);
  CarryOperator U240 (G4[40], P4[40], G3[40], P3[40], G3[32], P3[32]);
  CarryOperator U241 (G4[41], P4[41], G3[41], P3[41], G3[33], P3[33]);
  CarryOperator U242 (G4[42], P4[42], G3[42], P3[42], G3[34], P3[34]);
  CarryOperator U243 (G4[43], P4[43], G3[43], P3[43], G3[35], P3[35]);
  CarryOperator U244 (G4[44], P4[44], G3[44], P3[44], G3[36], P3[36]);
  CarryOperator U245 (G4[45], P4[45], G3[45], P3[45], G3[37], P3[37]);
  CarryOperator U246 (G4[46], P4[46], G3[46], P3[46], G3[38], P3[38]);
  CarryOperator U247 (G4[47], P4[47], G3[47], P3[47], G3[39], P3[39]);
  CarryOperator U248 (G4[48], P4[48], G3[48], P3[48], G3[40], P3[40]);
  CarryOperator U249 (G4[49], P4[49], G3[49], P3[49], G3[41], P3[41]);
  CarryOperator U250 (G4[50], P4[50], G3[50], P3[50], G3[42], P3[42]);
  CarryOperator U251 (G4[51], P4[51], G3[51], P3[51], G3[43], P3[43]);
  CarryOperator U252 (G4[52], P4[52], G3[52], P3[52], G3[44], P3[44]);
  CarryOperator U253 (G4[53], P4[53], G3[53], P3[53], G3[45], P3[45]);
  CarryOperator U254 (G4[54], P4[54], G3[54], P3[54], G3[46], P3[46]);
  CarryOperator U255 (G4[55], P4[55], G3[55], P3[55], G3[47], P3[47]);
  CarryOperator U256 (G4[56], P4[56], G3[56], P3[56], G3[48], P3[48]);
  CarryOperator U257 (G4[57], P4[57], G3[57], P3[57], G3[49], P3[49]);
  CarryOperator U258 (G4[58], P4[58], G3[58], P3[58], G3[50], P3[50]);
  CarryOperator U259 (G4[59], P4[59], G3[59], P3[59], G3[51], P3[51]);
  CarryOperator U260 (G4[60], P4[60], G3[60], P3[60], G3[52], P3[52]);
  CarryOperator U261 (G4[61], P4[61], G3[61], P3[61], G3[53], P3[53]);
  CarryOperator U262 (G4[62], P4[62], G3[62], P3[62], G3[54], P3[54]);
  CarryOperator U263 (G4[63], P4[63], G3[63], P3[63], G3[55], P3[55]);
  CarryOperator U264 (G4[64], P4[64], G3[64], P3[64], G3[56], P3[56]);
  CarryOperator U265 (G5[25], P5[25], G4[25], P4[25], G4[9], P4[9]);
  CarryOperator U266 (G5[26], P5[26], G4[26], P4[26], G4[10], P4[10]);
  CarryOperator U267 (G5[27], P5[27], G4[27], P4[27], G4[11], P4[11]);
  CarryOperator U268 (G5[28], P5[28], G4[28], P4[28], G4[12], P4[12]);
  CarryOperator U269 (G5[29], P5[29], G4[29], P4[29], G4[13], P4[13]);
  CarryOperator U270 (G5[30], P5[30], G4[30], P4[30], G4[14], P4[14]);
  CarryOperator U271 (G5[31], P5[31], G4[31], P4[31], G4[15], P4[15]);
  CarryOperator U272 (G5[32], P5[32], G4[32], P4[32], G4[16], P4[16]);
  CarryOperator U273 (G5[33], P5[33], G4[33], P4[33], G4[17], P4[17]);
  CarryOperator U274 (G5[34], P5[34], G4[34], P4[34], G4[18], P4[18]);
  CarryOperator U275 (G5[35], P5[35], G4[35], P4[35], G4[19], P4[19]);
  CarryOperator U276 (G5[36], P5[36], G4[36], P4[36], G4[20], P4[20]);
  CarryOperator U277 (G5[37], P5[37], G4[37], P4[37], G4[21], P4[21]);
  CarryOperator U278 (G5[38], P5[38], G4[38], P4[38], G4[22], P4[22]);
  CarryOperator U279 (G5[39], P5[39], G4[39], P4[39], G4[23], P4[23]);
  CarryOperator U280 (G5[40], P5[40], G4[40], P4[40], G4[24], P4[24]);
  CarryOperator U281 (G5[41], P5[41], G4[41], P4[41], G4[25], P4[25]);
  CarryOperator U282 (G5[42], P5[42], G4[42], P4[42], G4[26], P4[26]);
  CarryOperator U283 (G5[43], P5[43], G4[43], P4[43], G4[27], P4[27]);
  CarryOperator U284 (G5[44], P5[44], G4[44], P4[44], G4[28], P4[28]);
  CarryOperator U285 (G5[45], P5[45], G4[45], P4[45], G4[29], P4[29]);
  CarryOperator U286 (G5[46], P5[46], G4[46], P4[46], G4[30], P4[30]);
  CarryOperator U287 (G5[47], P5[47], G4[47], P4[47], G4[31], P4[31]);
  CarryOperator U288 (G5[48], P5[48], G4[48], P4[48], G4[32], P4[32]);
  CarryOperator U289 (G5[49], P5[49], G4[49], P4[49], G4[33], P4[33]);
  CarryOperator U290 (G5[50], P5[50], G4[50], P4[50], G4[34], P4[34]);
  CarryOperator U291 (G5[51], P5[51], G4[51], P4[51], G4[35], P4[35]);
  CarryOperator U292 (G5[52], P5[52], G4[52], P4[52], G4[36], P4[36]);
  CarryOperator U293 (G5[53], P5[53], G4[53], P4[53], G4[37], P4[37]);
  CarryOperator U294 (G5[54], P5[54], G4[54], P4[54], G4[38], P4[38]);
  CarryOperator U295 (G5[55], P5[55], G4[55], P4[55], G4[39], P4[39]);
  CarryOperator U296 (G5[56], P5[56], G4[56], P4[56], G4[40], P4[40]);
  CarryOperator U297 (G5[57], P5[57], G4[57], P4[57], G4[41], P4[41]);
  CarryOperator U298 (G5[58], P5[58], G4[58], P4[58], G4[42], P4[42]);
  CarryOperator U299 (G5[59], P5[59], G4[59], P4[59], G4[43], P4[43]);
  CarryOperator U300 (G5[60], P5[60], G4[60], P4[60], G4[44], P4[44]);
  CarryOperator U301 (G5[61], P5[61], G4[61], P4[61], G4[45], P4[45]);
  CarryOperator U302 (G5[62], P5[62], G4[62], P4[62], G4[46], P4[46]);
  CarryOperator U303 (G5[63], P5[63], G4[63], P4[63], G4[47], P4[47]);
  CarryOperator U304 (G5[64], P5[64], G4[64], P4[64], G4[48], P4[48]);
  CarryOperator U305 (G6[41], P6[41], G5[41], P5[41], G5[9], P5[9]);
  CarryOperator U306 (G6[42], P6[42], G5[42], P5[42], G5[10], P5[10]);
  CarryOperator U307 (G6[43], P6[43], G5[43], P5[43], G5[11], P5[11]);
  CarryOperator U308 (G6[44], P6[44], G5[44], P5[44], G5[12], P5[12]);
  CarryOperator U309 (G6[45], P6[45], G5[45], P5[45], G5[13], P5[13]);
  CarryOperator U310 (G6[46], P6[46], G5[46], P5[46], G5[14], P5[14]);
  CarryOperator U311 (G6[47], P6[47], G5[47], P5[47], G5[15], P5[15]);
  CarryOperator U312 (G6[48], P6[48], G5[48], P5[48], G5[16], P5[16]);
  CarryOperator U313 (G6[49], P6[49], G5[49], P5[49], G5[17], P5[17]);
  CarryOperator U314 (G6[50], P6[50], G5[50], P5[50], G5[18], P5[18]);
  CarryOperator U315 (G6[51], P6[51], G5[51], P5[51], G5[19], P5[19]);
  CarryOperator U316 (G6[52], P6[52], G5[52], P5[52], G5[20], P5[20]);
  CarryOperator U317 (G6[53], P6[53], G5[53], P5[53], G5[21], P5[21]);
  CarryOperator U318 (G6[54], P6[54], G5[54], P5[54], G5[22], P5[22]);
  CarryOperator U319 (G6[55], P6[55], G5[55], P5[55], G5[23], P5[23]);
  CarryOperator U320 (G6[56], P6[56], G5[56], P5[56], G5[24], P5[24]);
  CarryOperator U321 (G6[57], P6[57], G5[57], P5[57], G5[25], P5[25]);
  CarryOperator U322 (G6[58], P6[58], G5[58], P5[58], G5[26], P5[26]);
  CarryOperator U323 (G6[59], P6[59], G5[59], P5[59], G5[27], P5[27]);
  CarryOperator U324 (G6[60], P6[60], G5[60], P5[60], G5[28], P5[28]);
  CarryOperator U325 (G6[61], P6[61], G5[61], P5[61], G5[29], P5[29]);
  CarryOperator U326 (G6[62], P6[62], G5[62], P5[62], G5[30], P5[30]);
  CarryOperator U327 (G6[63], P6[63], G5[63], P5[63], G5[31], P5[31]);
  CarryOperator U328 (G6[64], P6[64], G5[64], P5[64], G5[32], P5[32]);
endmodule

module UBZero_9_9(O);
  output [9:9] O;
  assign O[9] = 0;
endmodule

module UBTC1CON66_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_32(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_33(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_34(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_35(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_36(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_37(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_38(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_39(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_40(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_41(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_42(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_43(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_44(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_45(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_46(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_47(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_48(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_49(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_50(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_51(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_52(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_53(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_54(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_55(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_56(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_57(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_58(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_59(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_60(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_61(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_62(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTCTCONV_65_63(O, I);
  output [66:63] O;
  input [65:63] I;
  assign O[63] = ~ I[63];
  assign O[64] = ~ I[64] ^ ( I[63] );
  assign O[65] = ~ I[65] ^ ( I[64] | I[63] );
  assign O[66] = ~ ( I[65] | I[64] | I[63] );
endmodule

module Multiplier_31_0_3000(P, IN1, IN2);

  output [63:0] P;
  input [31:0] IN1;
  input [31:0] IN2;
  wire [66:0] W;
  assign P[0] = W[0];
  assign P[1] = W[1];
  assign P[2] = W[2];
  assign P[3] = W[3];
  assign P[4] = W[4];
  assign P[5] = W[5];
  assign P[6] = W[6];
  assign P[7] = W[7];
  assign P[8] = W[8];
  assign P[9] = W[9];
  assign P[10] = W[10];
  assign P[11] = W[11];
  assign P[12] = W[12];
  assign P[13] = W[13];
  assign P[14] = W[14];
  assign P[15] = W[15];
  assign P[16] = W[16];
  assign P[17] = W[17];
  assign P[18] = W[18];
  assign P[19] = W[19];
  assign P[20] = W[20];
  assign P[21] = W[21];
  assign P[22] = W[22];
  assign P[23] = W[23];
  assign P[24] = W[24];
  assign P[25] = W[25];
  assign P[26] = W[26];
  assign P[27] = W[27];
  assign P[28] = W[28];
  assign P[29] = W[29];
  assign P[30] = W[30];
  assign P[31] = W[31];
  assign P[32] = W[32];
  assign P[33] = W[33];
  assign P[34] = W[34];
  assign P[35] = W[35];
  assign P[36] = W[36];
  assign P[37] = W[37];
  assign P[38] = W[38];
  assign P[39] = W[39];
  assign P[40] = W[40];
  assign P[41] = W[41];
  assign P[42] = W[42];
  assign P[43] = W[43];
  assign P[44] = W[44];
  assign P[45] = W[45];
  assign P[46] = W[46];
  assign P[47] = W[47];
  assign P[48] = W[48];
  assign P[49] = W[49];
  assign P[50] = W[50];
  assign P[51] = W[51];
  assign P[52] = W[52];
  assign P[53] = W[53];
  assign P[54] = W[54];
  assign P[55] = W[55];
  assign P[56] = W[56];
  assign P[57] = W[57];
  assign P[58] = W[58];
  assign P[59] = W[59];
  assign P[60] = W[60];
  assign P[61] = W[61];
  assign P[62] = W[62];
  assign P[63] = W[63];
  MultTC_STD_WAL_KS000 U0 (W, IN1, IN2);
endmodule

module CSA_32_0_32_1_33_000 (C, S, X, Y, Z);
  output [33:2] C;
  output [33:0] S;
  input [32:0] X;
  input [32:1] Y;
  input [33:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_32_2 U2 (C[33:3], S[32:2], Z[32:2], Y[32:2], X[32:2]);
  UB1DCON_33 U3 (S[33], Z[33]);
endmodule

module CSA_33_0_33_2_36_000 (C, S, X, Y, Z);
  output [34:3] C;
  output [36:0] S;
  input [33:0] X;
  input [33:2] Y;
  input [36:3] Z;
  UBCON_1_0 U0 (S[1:0], X[1:0]);
  UBHA_2 U1 (C[3], S[2], Y[2], X[2]);
  PureCSA_33_3 U2 (C[34:4], S[33:3], Z[33:3], Y[33:3], X[33:3]);
  UBCON_36_34 U3 (S[36:34], Z[36:34]);
endmodule

module CSA_34_3_35_4_36_000 (C, S, X, Y, Z);
  output [36:5] C;
  output [36:3] S;
  input [34:3] X;
  input [35:4] Y;
  input [36:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_34_5 U2 (C[35:6], S[34:5], Z[34:5], Y[34:5], X[34:5]);
  UBHA_35 U3 (C[36], S[35], Z[35], Y[35]);
  UB1DCON_36 U4 (S[36], Z[36]);
endmodule

module CSA_36_0_34_3_39_000 (C, S, X, Y, Z);
  output [37:4] C;
  output [39:0] S;
  input [36:0] X;
  input [34:3] Y;
  input [39:5] Z;
  UBCON_2_0 U0 (S[2:0], X[2:0]);
  PureCSHA_4_3 U1 (C[5:4], S[4:3], Y[4:3], X[4:3]);
  PureCSA_34_5 U2 (C[35:6], S[34:5], Z[34:5], Y[34:5], X[34:5]);
  PureCSHA_36_35 U3 (C[37:36], S[36:35], Z[36:35], X[36:35]);
  UBCON_39_37 U4 (S[39:37], Z[39:37]);
endmodule

module CSA_36_5_39_6_39_000 (C, S, X, Y, Z);
  output [40:7] C;
  output [39:5] S;
  input [36:5] X;
  input [39:6] Y;
  input [39:8] Z;
  UB1DCON_5 U0 (S[5], X[5]);
  PureCSHA_7_6 U1 (C[8:7], S[7:6], Y[7:6], X[7:6]);
  PureCSA_36_8 U2 (C[37:9], S[36:8], Z[36:8], Y[36:8], X[36:8]);
  PureCSHA_39_37 U3 (C[40:38], S[39:37], Z[39:37], Y[39:37]);
endmodule

module CSA_37_6_38_7_39_000 (C, S, X, Y, Z);
  output [39:8] C;
  output [39:6] S;
  input [37:6] X;
  input [38:7] Y;
  input [39:8] Z;
  UB1DCON_6 U0 (S[6], X[6]);
  UBHA_7 U1 (C[8], S[7], Y[7], X[7]);
  PureCSA_37_8 U2 (C[38:9], S[37:8], Z[37:8], Y[37:8], X[37:8]);
  UBHA_38 U3 (C[39], S[38], Z[38], Y[38]);
  UB1DCON_39 U4 (S[39], Z[39]);
endmodule

module CSA_39_0_37_4_43_000 (C, S, X, Y, Z);
  output [40:5] C;
  output [43:0] S;
  input [39:0] X;
  input [37:4] Y;
  input [43:7] Z;
  UBCON_3_0 U0 (S[3:0], X[3:0]);
  PureCSHA_6_4 U1 (C[7:5], S[6:4], Y[6:4], X[6:4]);
  PureCSA_37_7 U2 (C[38:8], S[37:7], Z[37:7], Y[37:7], X[37:7]);
  PureCSHA_39_38 U3 (C[40:39], S[39:38], Z[39:38], X[39:38]);
  UBCON_43_40 U4 (S[43:40], Z[43:40]);
endmodule

module CSA_40_7_43_9_43_000 (C, S, X, Y, Z);
  output [44:10] C;
  output [43:7] S;
  input [40:7] X;
  input [43:9] Y;
  input [43:12] Z;
  UBCON_8_7 U0 (S[8:7], X[8:7]);
  PureCSHA_11_9 U1 (C[12:10], S[11:9], Y[11:9], X[11:9]);
  PureCSA_40_12 U2 (C[41:13], S[40:12], Z[40:12], Y[40:12], X[40:12]);
  PureCSHA_43_41 U3 (C[44:42], S[43:41], Z[43:41], Y[43:41]);
endmodule

module CSA_40_9_41_10_42000 (C, S, X, Y, Z);
  output [42:11] C;
  output [42:9] S;
  input [40:9] X;
  input [41:10] Y;
  input [42:11] Z;
  UB1DCON_9 U0 (S[9], X[9]);
  UBHA_10 U1 (C[11], S[10], Y[10], X[10]);
  PureCSA_40_11 U2 (C[41:12], S[40:11], Z[40:11], Y[40:11], X[40:11]);
  UBHA_41 U3 (C[42], S[41], Z[41], Y[41]);
  UB1DCON_42 U4 (S[42], Z[42]);
endmodule

module CSA_42_9_42_11_43000 (C, S, X, Y, Z);
  output [43:12] C;
  output [43:9] S;
  input [42:9] X;
  input [42:11] Y;
  input [43:12] Z;
  UBCON_10_9 U0 (S[10:9], X[10:9]);
  UBHA_11 U1 (C[12], S[11], Y[11], X[11]);
  PureCSA_42_12 U2 (C[43:13], S[42:12], Z[42:12], Y[42:12], X[42:12]);
  UB1DCON_43 U3 (S[43], Z[43]);
endmodule

module CSA_43_0_40_5_49_000 (C, S, X, Y, Z);
  output [44:6] C;
  output [49:0] S;
  input [43:0] X;
  input [40:5] Y;
  input [49:10] Z;
  UBCON_4_0 U0 (S[4:0], X[4:0]);
  PureCSHA_9_5 U1 (C[10:6], S[9:5], Y[9:5], X[9:5]);
  PureCSA_40_10 U2 (C[41:11], S[40:10], Z[40:10], Y[40:10], X[40:10]);
  PureCSHA_43_41 U3 (C[44:42], S[43:41], Z[43:41], X[43:41]);
  UBCON_49_44 U4 (S[49:44], Z[49:44]);
endmodule

module CSA_44_10_49_13_4000 (C, S, X, Y, Z);
  output [48:14] C;
  output [49:10] S;
  input [44:10] X;
  input [49:13] Y;
  input [47:16] Z;
  UBCON_12_10 U0 (S[12:10], X[12:10]);
  PureCSHA_15_13 U1 (C[16:14], S[15:13], Y[15:13], X[15:13]);
  PureCSA_44_16 U2 (C[45:17], S[44:16], Z[44:16], Y[44:16], X[44:16]);
  PureCSHA_47_45 U3 (C[48:46], S[47:45], Y[47:45], Z[47:45]);
  UBCON_49_48 U4 (S[49:48], Y[49:48]);
endmodule

module CSA_44_13_45_14_4000 (C, S, X, Y, Z);
  output [46:15] C;
  output [46:13] S;
  input [44:13] X;
  input [45:14] Y;
  input [46:15] Z;
  UB1DCON_13 U0 (S[13], X[13]);
  UBHA_14 U1 (C[15], S[14], Y[14], X[14]);
  PureCSA_44_15 U2 (C[45:16], S[44:15], Z[44:15], Y[44:15], X[44:15]);
  UBHA_45 U3 (C[46], S[45], Z[45], Y[45]);
  UB1DCON_46 U4 (S[46], Z[46]);
endmodule

module CSA_46_13_46_15_4000 (C, S, X, Y, Z);
  output [47:16] C;
  output [49:13] S;
  input [46:13] X;
  input [46:15] Y;
  input [49:16] Z;
  UBCON_14_13 U0 (S[14:13], X[14:13]);
  UBHA_15 U1 (C[16], S[15], Y[15], X[15]);
  PureCSA_46_16 U2 (C[47:17], S[46:16], Z[46:16], Y[46:16], X[46:16]);
  UBCON_49_47 U3 (S[49:47], Z[49:47]);
endmodule

module CSA_47_16_48_17_4000 (C, S, X, Y, Z);
  output [49:18] C;
  output [49:16] S;
  input [47:16] X;
  input [48:17] Y;
  input [49:18] Z;
  UB1DCON_16 U0 (S[16], X[16]);
  UBHA_17 U1 (C[18], S[17], Y[17], X[17]);
  PureCSA_47_18 U2 (C[48:19], S[47:18], Z[47:18], Y[47:18], X[47:18]);
  UBHA_48 U3 (C[49], S[48], Z[48], Y[48]);
  UB1DCON_49 U4 (S[49], Z[49]);
endmodule

module CSA_48_14_58_18_5000 (C, S, X, Y, Z);
  output [55:19] C;
  output [58:14] S;
  input [48:14] X;
  input [58:18] Y;
  input [54:21] Z;
  UBCON_17_14 U0 (S[17:14], X[17:14]);
  PureCSHA_20_18 U1 (C[21:19], S[20:18], Y[20:18], X[20:18]);
  PureCSA_48_21 U2 (C[49:22], S[48:21], Z[48:21], Y[48:21], X[48:21]);
  PureCSHA_54_49 U3 (C[55:50], S[54:49], Y[54:49], Z[54:49]);
  UBCON_58_55 U4 (S[58:55], Y[58:55]);
endmodule

module CSA_49_0_44_6_58_000 (C, S, X, Y, Z);
  output [50:7] C;
  output [58:0] S;
  input [49:0] X;
  input [44:6] Y;
  input [58:14] Z;
  UBCON_5_0 U0 (S[5:0], X[5:0]);
  PureCSHA_13_6 U1 (C[14:7], S[13:6], Y[13:6], X[13:6]);
  PureCSA_44_14 U2 (C[45:15], S[44:14], Z[44:14], Y[44:14], X[44:14]);
  PureCSHA_49_45 U3 (C[50:46], S[49:45], Z[49:45], X[49:45]);
  UBCON_58_50 U4 (S[58:50], Z[58:50]);
endmodule

module CSA_49_18_52_19_5000 (C, S, X, Y, Z);
  output [53:20] C;
  output [52:18] S;
  input [49:18] X;
  input [52:19] Y;
  input [52:21] Z;
  UB1DCON_18 U0 (S[18], X[18]);
  PureCSHA_20_19 U1 (C[21:20], S[20:19], Y[20:19], X[20:19]);
  PureCSA_49_21 U2 (C[50:22], S[49:21], Z[49:21], Y[49:21], X[49:21]);
  PureCSHA_52_50 U3 (C[53:51], S[52:50], Z[52:50], Y[52:50]);
endmodule

module CSA_50_19_51_20_5000 (C, S, X, Y, Z);
  output [52:21] C;
  output [52:19] S;
  input [50:19] X;
  input [51:20] Y;
  input [52:21] Z;
  UB1DCON_19 U0 (S[19], X[19]);
  UBHA_20 U1 (C[21], S[20], Y[20], X[20]);
  PureCSA_50_21 U2 (C[51:22], S[50:21], Z[50:21], Y[50:21], X[50:21]);
  UBHA_51 U3 (C[52], S[51], Z[51], Y[51]);
  UB1DCON_52 U4 (S[52], Z[52]);
endmodule

module CSA_52_18_53_20_5000 (C, S, X, Y, Z);
  output [54:21] C;
  output [58:18] S;
  input [52:18] X;
  input [53:20] Y;
  input [58:22] Z;
  UBCON_19_18 U0 (S[19:18], X[19:18]);
  PureCSHA_21_20 U1 (C[22:21], S[21:20], Y[21:20], X[21:20]);
  PureCSA_52_22 U2 (C[53:23], S[52:22], Z[52:22], Y[52:22], X[52:22]);
  UBHA_53 U3 (C[54], S[53], Z[53], Y[53]);
  UBCON_58_54 U4 (S[58:54], Z[58:54]);
endmodule

module CSA_53_22_54_23_5000 (C, S, X, Y, Z);
  output [55:24] C;
  output [55:22] S;
  input [53:22] X;
  input [54:23] Y;
  input [55:24] Z;
  UB1DCON_22 U0 (S[22], X[22]);
  UBHA_23 U1 (C[24], S[23], Y[23], X[23]);
  PureCSA_53_24 U2 (C[54:25], S[53:24], Z[53:24], Y[53:24], X[53:24]);
  UBHA_54 U3 (C[55], S[54], Z[54], Y[54]);
  UB1DCON_55 U4 (S[55], Z[55]);
endmodule

module CSA_55_19_62_25_6000 (C, S, X, Y, Z);
  output [63:26] C;
  output [63:19] S;
  input [55:19] X;
  input [62:25] Y;
  input [63:29] Z;
  UBCON_24_19 U0 (S[24:19], X[24:19]);
  PureCSHA_28_25 U1 (C[29:26], S[28:25], Y[28:25], X[28:25]);
  PureCSA_55_29 U2 (C[56:30], S[55:29], Z[55:29], Y[55:29], X[55:29]);
  PureCSHA_62_56 U3 (C[63:57], S[62:56], Z[62:56], Y[62:56]);
  UB1DCON_63 U4 (S[63], Z[63]);
endmodule

module CSA_55_22_55_24_5000 (C, S, X, Y, Z);
  output [56:25] C;
  output [58:22] S;
  input [55:22] X;
  input [55:24] Y;
  input [58:25] Z;
  UBCON_23_22 U0 (S[23:22], X[23:22]);
  UBHA_24 U1 (C[25], S[24], Y[24], X[24]);
  PureCSA_55_25 U2 (C[56:26], S[55:25], Z[55:25], Y[55:25], X[55:25]);
  UBCON_58_56 U3 (S[58:56], Z[58:56]);
endmodule

module CSA_56_25_57_26_5000 (C, S, X, Y, Z);
  output [58:27] C;
  output [58:25] S;
  input [56:25] X;
  input [57:26] Y;
  input [58:27] Z;
  UB1DCON_25 U0 (S[25], X[25]);
  UBHA_26 U1 (C[27], S[26], Y[26], X[26]);
  PureCSA_56_27 U2 (C[57:28], S[56:27], Z[56:27], Y[56:27], X[56:27]);
  UBHA_57 U3 (C[58], S[57], Z[57], Y[57]);
  UB1DCON_58 U4 (S[58], Z[58]);
endmodule

module CSA_56_25_61_27_6000 (C, S, X, Y, Z);
  output [62:28] C;
  output [62:25] S;
  input [56:25] X;
  input [61:27] Y;
  input [62:29] Z;
  UBCON_26_25 U0 (S[26:25], X[26:25]);
  PureCSHA_28_27 U1 (C[29:28], S[28:27], Y[28:27], X[28:27]);
  PureCSA_56_29 U2 (C[57:30], S[56:29], Z[56:29], Y[56:29], X[56:29]);
  PureCSHA_61_57 U3 (C[62:58], S[61:57], Z[61:57], Y[61:57]);
  UB1DCON_62 U4 (S[62], Z[62]);
endmodule

module CSA_58_0_50_7_63_000 (C, S, X, Y, Z);
  output [59:8] C;
  output [63:0] S;
  input [58:0] X;
  input [50:7] Y;
  input [63:19] Z;
  UBCON_6_0 U0 (S[6:0], X[6:0]);
  PureCSHA_18_7 U1 (C[19:8], S[18:7], Y[18:7], X[18:7]);
  PureCSA_50_19 U2 (C[51:20], S[50:19], Z[50:19], Y[50:19], X[50:19]);
  PureCSHA_58_51 U3 (C[59:52], S[58:51], Z[58:51], X[58:51]);
  UBCON_63_59 U4 (S[63:59], Z[63:59]);
endmodule

module CSA_58_27_61_28_6000 (C, S, X, Y, Z);
  output [62:29] C;
  output [61:27] S;
  input [58:27] X;
  input [61:28] Y;
  input [61:30] Z;
  UB1DCON_27 U0 (S[27], X[27]);
  PureCSHA_29_28 U1 (C[30:29], S[29:28], Y[29:28], X[29:28]);
  PureCSA_58_30 U2 (C[59:31], S[58:30], Z[58:30], Y[58:30], X[58:30]);
  PureCSHA_61_59 U3 (C[62:60], S[61:59], Z[61:59], Y[61:59]);
endmodule

module CSA_59_28_60_29_6000 (C, S, X, Y, Z);
  output [61:30] C;
  output [61:28] S;
  input [59:28] X;
  input [60:29] Y;
  input [61:30] Z;
  UB1DCON_28 U0 (S[28], X[28]);
  UBHA_29 U1 (C[30], S[29], Y[29], X[29]);
  PureCSA_59_30 U2 (C[60:31], S[59:30], Z[59:30], Y[59:30], X[59:30]);
  UBHA_60 U3 (C[61], S[60], Z[60], Y[60]);
  UB1DCON_61 U4 (S[61], Z[61]);
endmodule

module CSA_62_25_62_28_6000 (C, S, X, Y, Z);
  output [63:29] C;
  output [62:25] S;
  input [62:25] X;
  input [62:28] Y;
  input [62:31] Z;
  UBCON_27_25 U0 (S[27:25], X[27:25]);
  PureCSHA_30_28 U1 (C[31:29], S[30:28], Y[30:28], X[30:28]);
  PureCSA_62_31 U2 (C[63:32], S[62:31], Z[62:31], Y[62:31], X[62:31]);
endmodule

module CSA_63_0_59_8_63_000 (C, S, X, Y, Z);
  output [64:9] C;
  output [63:0] S;
  input [63:0] X;
  input [59:8] Y;
  input [63:26] Z;
  UBCON_7_0 U0 (S[7:0], X[7:0]);
  PureCSHA_25_8 U1 (C[26:9], S[25:8], Y[25:8], X[25:8]);
  PureCSA_59_26 U2 (C[60:27], S[59:26], Z[59:26], Y[59:26], X[59:26]);
  PureCSHA_63_60 U3 (C[64:61], S[63:60], Z[63:60], X[63:60]);
endmodule

module MultTC_STD_WAL_KS000 (P, IN1, IN2);

  output [66:0] P;
  input [31:0] IN1;
  input [31:0] IN2;
  wire [32:0] PP0;
  wire [32:1] PP1;
  wire [41:10] PP10;
  wire [42:11] PP11;
  wire [43:12] PP12;
  wire [44:13] PP13;
  wire [45:14] PP14;
  wire [46:15] PP15;
  wire [47:16] PP16;
  wire [48:17] PP17;
  wire [49:18] PP18;
  wire [50:19] PP19;
  wire [33:2] PP2;
  wire [51:20] PP20;
  wire [52:21] PP21;
  wire [53:22] PP22;
  wire [54:23] PP23;
  wire [55:24] PP24;
  wire [56:25] PP25;
  wire [57:26] PP26;
  wire [58:27] PP27;
  wire [59:28] PP28;
  wire [60:29] PP29;
  wire [34:3] PP3;
  wire [61:30] PP30;
  wire [62:31] PP31;
  wire [35:4] PP4;
  wire [36:5] PP5;
  wire [37:6] PP6;
  wire [38:7] PP7;
  wire [39:8] PP8;
  wire [40:9] PP9;
  wire [65:0] P_UB;
  wire [64:9] S1;
  wire [63:0] S2;

  TCPPG_31_0_31_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, IN1, IN2);
  WLCTR_32_0_32_1_3000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31);

  UBKSA_64_9_63_0 U2 (P_UB, S1, S2);
  UBTCCONV63_65_0 U3 (P, P_UB);
endmodule

module NUBUBCON_61_31 (O, I);
  output [61:31] O;
  input [61:31] I;
  NUBUB1CON_31 U0 (O[31], I[31]);
  NUBUB1CON_32 U1 (O[32], I[32]);
  NUBUB1CON_33 U2 (O[33], I[33]);
  NUBUB1CON_34 U3 (O[34], I[34]);
  NUBUB1CON_35 U4 (O[35], I[35]);
  NUBUB1CON_36 U5 (O[36], I[36]);
  NUBUB1CON_37 U6 (O[37], I[37]);
  NUBUB1CON_38 U7 (O[38], I[38]);
  NUBUB1CON_39 U8 (O[39], I[39]);
  NUBUB1CON_40 U9 (O[40], I[40]);
  NUBUB1CON_41 U10 (O[41], I[41]);
  NUBUB1CON_42 U11 (O[42], I[42]);
  NUBUB1CON_43 U12 (O[43], I[43]);
  NUBUB1CON_44 U13 (O[44], I[44]);
  NUBUB1CON_45 U14 (O[45], I[45]);
  NUBUB1CON_46 U15 (O[46], I[46]);
  NUBUB1CON_47 U16 (O[47], I[47]);
  NUBUB1CON_48 U17 (O[48], I[48]);
  NUBUB1CON_49 U18 (O[49], I[49]);
  NUBUB1CON_50 U19 (O[50], I[50]);
  NUBUB1CON_51 U20 (O[51], I[51]);
  NUBUB1CON_52 U21 (O[52], I[52]);
  NUBUB1CON_53 U22 (O[53], I[53]);
  NUBUB1CON_54 U23 (O[54], I[54]);
  NUBUB1CON_55 U24 (O[55], I[55]);
  NUBUB1CON_56 U25 (O[56], I[56]);
  NUBUB1CON_57 U26 (O[57], I[57]);
  NUBUB1CON_58 U27 (O[58], I[58]);
  NUBUB1CON_59 U28 (O[59], I[59]);
  NUBUB1CON_60 U29 (O[60], I[60]);
  NUBUB1CON_61 U30 (O[61], I[61]);
endmodule

module PureCSA_32_2 (C, S, X, Y, Z);
  output [33:3] C;
  output [32:2] S;
  input [32:2] X;
  input [32:2] Y;
  input [32:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U4 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U5 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U6 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U7 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U8 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U9 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U10 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U11 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U12 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U13 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U14 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U15 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U16 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U17 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U18 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U19 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U20 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U21 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U22 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U23 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U24 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U25 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U26 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U27 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U28 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U29 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U30 (C[33], S[32], X[32], Y[32], Z[32]);
endmodule

module PureCSA_33_3 (C, S, X, Y, Z);
  output [34:4] C;
  output [33:3] S;
  input [33:3] X;
  input [33:3] Y;
  input [33:3] Z;
  UBFA_3 U0 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U1 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U2 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U3 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U4 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U5 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U6 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U7 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U8 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U9 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U10 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U11 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U12 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U13 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U14 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U15 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U16 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U17 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U18 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U19 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U20 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U21 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U22 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U23 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U24 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U25 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U26 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U27 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U28 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U29 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U30 (C[34], S[33], X[33], Y[33], Z[33]);
endmodule

module PureCSA_34_5 (C, S, X, Y, Z);
  output [35:6] C;
  output [34:5] S;
  input [34:5] X;
  input [34:5] Y;
  input [34:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U7 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U8 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U9 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U10 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U11 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U12 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U13 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U14 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U15 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U16 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U17 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U18 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U19 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U20 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U21 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U22 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U23 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U24 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U25 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U26 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U27 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U28 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U29 (C[35], S[34], X[34], Y[34], Z[34]);
endmodule

module PureCSA_36_8 (C, S, X, Y, Z);
  output [37:9] C;
  output [36:8] S;
  input [36:8] X;
  input [36:8] Y;
  input [36:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U11 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U12 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U13 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U14 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U15 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U16 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U17 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U18 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U19 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U20 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U21 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U22 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U23 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U24 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U25 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U26 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U27 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U28 (C[37], S[36], X[36], Y[36], Z[36]);
endmodule

module PureCSA_37_7 (C, S, X, Y, Z);
  output [38:8] C;
  output [37:7] S;
  input [37:7] X;
  input [37:7] Y;
  input [37:7] Z;
  UBFA_7 U0 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U1 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U2 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U3 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U4 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U5 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U6 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U7 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U8 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U9 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U10 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U11 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U12 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U13 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U14 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U15 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U16 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U17 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U18 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U19 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U20 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U21 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U22 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U23 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U24 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U25 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U26 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U27 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U28 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U29 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U30 (C[38], S[37], X[37], Y[37], Z[37]);
endmodule

module PureCSA_37_8 (C, S, X, Y, Z);
  output [38:9] C;
  output [37:8] S;
  input [37:8] X;
  input [37:8] Y;
  input [37:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U11 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U12 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U13 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U14 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U15 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U16 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U17 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U18 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U19 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U20 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U21 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U22 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U23 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U24 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U25 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U26 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U27 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U28 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U29 (C[38], S[37], X[37], Y[37], Z[37]);
endmodule

module PureCSA_40_10 (C, S, X, Y, Z);
  output [41:11] C;
  output [40:10] S;
  input [40:10] X;
  input [40:10] Y;
  input [40:10] Z;
  UBFA_10 U0 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U1 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U2 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U3 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U4 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U5 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U6 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U7 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U8 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U9 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U10 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U11 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U12 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U13 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U14 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U15 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U16 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U17 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U18 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U19 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U20 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U21 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U22 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U23 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U24 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U25 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U26 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U27 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U28 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U29 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U30 (C[41], S[40], X[40], Y[40], Z[40]);
endmodule

module PureCSA_40_11 (C, S, X, Y, Z);
  output [41:12] C;
  output [40:11] S;
  input [40:11] X;
  input [40:11] Y;
  input [40:11] Z;
  UBFA_11 U0 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U1 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U2 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U3 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U4 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U5 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U6 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U7 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U8 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U9 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U10 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U11 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U12 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U13 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U14 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U15 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U16 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U17 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U18 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U19 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U20 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U21 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U22 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U23 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U24 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U25 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U26 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U27 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U28 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U29 (C[41], S[40], X[40], Y[40], Z[40]);
endmodule

module PureCSA_40_12 (C, S, X, Y, Z);
  output [41:13] C;
  output [40:12] S;
  input [40:12] X;
  input [40:12] Y;
  input [40:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U10 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U11 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U12 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U13 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U14 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U15 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U16 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U17 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U18 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U19 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U20 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U21 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U22 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U23 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U24 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U25 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U26 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U27 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U28 (C[41], S[40], X[40], Y[40], Z[40]);
endmodule

module PureCSA_42_12 (C, S, X, Y, Z);
  output [43:13] C;
  output [42:12] S;
  input [42:12] X;
  input [42:12] Y;
  input [42:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U10 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U11 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U12 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U13 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U14 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U15 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U16 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U17 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U18 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U19 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U20 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U21 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U22 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U23 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U24 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U25 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U26 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U27 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U28 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U29 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U30 (C[43], S[42], X[42], Y[42], Z[42]);
endmodule

module PureCSA_44_14 (C, S, X, Y, Z);
  output [45:15] C;
  output [44:14] S;
  input [44:14] X;
  input [44:14] Y;
  input [44:14] Z;
  UBFA_14 U0 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U1 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U2 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U3 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U4 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U5 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U6 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U7 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U8 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U9 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U10 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U11 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U12 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U13 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U14 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U15 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U16 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U17 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U18 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U19 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U20 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U21 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U22 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U23 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U24 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U25 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U26 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U27 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U28 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U29 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U30 (C[45], S[44], X[44], Y[44], Z[44]);
endmodule

module PureCSA_44_15 (C, S, X, Y, Z);
  output [45:16] C;
  output [44:15] S;
  input [44:15] X;
  input [44:15] Y;
  input [44:15] Z;
  UBFA_15 U0 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U1 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U2 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U3 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U4 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U5 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U6 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U7 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U8 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U9 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U10 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U11 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U12 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U13 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U14 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U15 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U16 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U17 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U18 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U19 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U20 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U21 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U22 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U23 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U24 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U25 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U26 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U27 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U28 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U29 (C[45], S[44], X[44], Y[44], Z[44]);
endmodule

module PureCSA_44_16 (C, S, X, Y, Z);
  output [45:17] C;
  output [44:16] S;
  input [44:16] X;
  input [44:16] Y;
  input [44:16] Z;
  UBFA_16 U0 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U1 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U2 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U3 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U4 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U5 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U6 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U7 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U8 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U9 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U10 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U11 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U12 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U13 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U14 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U15 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U16 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U17 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U18 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U19 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U20 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U21 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U22 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U23 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U24 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U25 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U26 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U27 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U28 (C[45], S[44], X[44], Y[44], Z[44]);
endmodule

module PureCSA_46_16 (C, S, X, Y, Z);
  output [47:17] C;
  output [46:16] S;
  input [46:16] X;
  input [46:16] Y;
  input [46:16] Z;
  UBFA_16 U0 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U1 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U2 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U3 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U4 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U5 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U6 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U7 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U8 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U9 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U10 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U11 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U12 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U13 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U14 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U15 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U16 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U17 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U18 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U19 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U20 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U21 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U22 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U23 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U24 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U25 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U26 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U27 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U28 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U29 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U30 (C[47], S[46], X[46], Y[46], Z[46]);
endmodule

module PureCSA_47_18 (C, S, X, Y, Z);
  output [48:19] C;
  output [47:18] S;
  input [47:18] X;
  input [47:18] Y;
  input [47:18] Z;
  UBFA_18 U0 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U1 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U2 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U3 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U4 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U5 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U6 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U7 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U8 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U9 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U10 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U11 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U12 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U13 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U14 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U15 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U16 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U17 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U18 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U19 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U20 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U21 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U22 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U23 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U24 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U25 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U26 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U27 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U28 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U29 (C[48], S[47], X[47], Y[47], Z[47]);
endmodule

module PureCSA_48_21 (C, S, X, Y, Z);
  output [49:22] C;
  output [48:21] S;
  input [48:21] X;
  input [48:21] Y;
  input [48:21] Z;
  UBFA_21 U0 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U1 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U2 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U3 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U4 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U5 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U6 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U7 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U8 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U9 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U10 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U11 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U12 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U13 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U14 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U15 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U16 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U17 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U18 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U19 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U20 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U21 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U22 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U23 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U24 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U25 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U26 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U27 (C[49], S[48], X[48], Y[48], Z[48]);
endmodule

module PureCSA_49_21 (C, S, X, Y, Z);
  output [50:22] C;
  output [49:21] S;
  input [49:21] X;
  input [49:21] Y;
  input [49:21] Z;
  UBFA_21 U0 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U1 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U2 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U3 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U4 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U5 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U6 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U7 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U8 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U9 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U10 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U11 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U12 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U13 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U14 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U15 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U16 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U17 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U18 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U19 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U20 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U21 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U22 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U23 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U24 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U25 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U26 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U27 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U28 (C[50], S[49], X[49], Y[49], Z[49]);
endmodule

module PureCSA_50_19 (C, S, X, Y, Z);
  output [51:20] C;
  output [50:19] S;
  input [50:19] X;
  input [50:19] Y;
  input [50:19] Z;
  UBFA_19 U0 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U1 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U2 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U3 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U4 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U5 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U6 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U7 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U8 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U9 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U10 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U11 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U12 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U13 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U14 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U15 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U16 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U17 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U18 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U19 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U20 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U21 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U22 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U23 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U24 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U25 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U26 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U27 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U28 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U29 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U30 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U31 (C[51], S[50], X[50], Y[50], Z[50]);
endmodule

module PureCSA_50_21 (C, S, X, Y, Z);
  output [51:22] C;
  output [50:21] S;
  input [50:21] X;
  input [50:21] Y;
  input [50:21] Z;
  UBFA_21 U0 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U1 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U2 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U3 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U4 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U5 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U6 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U7 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U8 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U9 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U10 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U11 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U12 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U13 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U14 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U15 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U16 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U17 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U18 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U19 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U20 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U21 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U22 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U23 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U24 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U25 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U26 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U27 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U28 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U29 (C[51], S[50], X[50], Y[50], Z[50]);
endmodule

module PureCSA_52_22 (C, S, X, Y, Z);
  output [53:23] C;
  output [52:22] S;
  input [52:22] X;
  input [52:22] Y;
  input [52:22] Z;
  UBFA_22 U0 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U1 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U2 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U3 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U4 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U5 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U6 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U7 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U8 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U9 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U10 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U11 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U12 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U13 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U14 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U15 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U16 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U17 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U18 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U19 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U20 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U21 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U22 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U23 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U24 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U25 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U26 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U27 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U28 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U29 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U30 (C[53], S[52], X[52], Y[52], Z[52]);
endmodule

module PureCSA_53_24 (C, S, X, Y, Z);
  output [54:25] C;
  output [53:24] S;
  input [53:24] X;
  input [53:24] Y;
  input [53:24] Z;
  UBFA_24 U0 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U1 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U2 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U3 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U4 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U5 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U6 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U7 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U8 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U9 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U10 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U11 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U12 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U13 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U14 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U15 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U16 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U17 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U18 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U19 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U20 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U21 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U22 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U23 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U24 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U25 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U26 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U27 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U28 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U29 (C[54], S[53], X[53], Y[53], Z[53]);
endmodule

module PureCSA_55_25 (C, S, X, Y, Z);
  output [56:26] C;
  output [55:25] S;
  input [55:25] X;
  input [55:25] Y;
  input [55:25] Z;
  UBFA_25 U0 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U1 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U2 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U3 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U4 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U5 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U6 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U7 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U8 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U9 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U10 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U11 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U12 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U13 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U14 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U15 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U16 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U17 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U18 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U19 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U20 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U21 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U22 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U23 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U24 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U25 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U26 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U27 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U28 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U29 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U30 (C[56], S[55], X[55], Y[55], Z[55]);
endmodule

module PureCSA_55_29 (C, S, X, Y, Z);
  output [56:30] C;
  output [55:29] S;
  input [55:29] X;
  input [55:29] Y;
  input [55:29] Z;
  UBFA_29 U0 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U1 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U2 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U3 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U4 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U5 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U6 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U7 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U8 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U9 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U10 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U11 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U12 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U13 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U14 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U15 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U16 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U17 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U18 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U19 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U20 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U21 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U22 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U23 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U24 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U25 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U26 (C[56], S[55], X[55], Y[55], Z[55]);
endmodule

module PureCSA_56_27 (C, S, X, Y, Z);
  output [57:28] C;
  output [56:27] S;
  input [56:27] X;
  input [56:27] Y;
  input [56:27] Z;
  UBFA_27 U0 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U1 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U2 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U3 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U4 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U5 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U6 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U7 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U8 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U9 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U10 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U11 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U12 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U13 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U14 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U15 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U16 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U17 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U18 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U19 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U20 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U21 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U22 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U23 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U24 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U25 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U26 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U27 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U28 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U29 (C[57], S[56], X[56], Y[56], Z[56]);
endmodule

module PureCSA_56_29 (C, S, X, Y, Z);
  output [57:30] C;
  output [56:29] S;
  input [56:29] X;
  input [56:29] Y;
  input [56:29] Z;
  UBFA_29 U0 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U1 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U2 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U3 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U4 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U5 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U6 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U7 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U8 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U9 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U10 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U11 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U12 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U13 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U14 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U15 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U16 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U17 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U18 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U19 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U20 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U21 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U22 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U23 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U24 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U25 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U26 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U27 (C[57], S[56], X[56], Y[56], Z[56]);
endmodule

module PureCSA_58_30 (C, S, X, Y, Z);
  output [59:31] C;
  output [58:30] S;
  input [58:30] X;
  input [58:30] Y;
  input [58:30] Z;
  UBFA_30 U0 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U1 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U2 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U3 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U4 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U5 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U6 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U7 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U8 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U9 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U10 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U11 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U12 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U13 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U14 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U15 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U16 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U17 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U18 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U19 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U20 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U21 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U22 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U23 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U24 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U25 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U26 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U27 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U28 (C[59], S[58], X[58], Y[58], Z[58]);
endmodule

module PureCSA_59_26 (C, S, X, Y, Z);
  output [60:27] C;
  output [59:26] S;
  input [59:26] X;
  input [59:26] Y;
  input [59:26] Z;
  UBFA_26 U0 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U1 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U2 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U3 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U4 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U5 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U6 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U7 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U8 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U9 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U10 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U11 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U12 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U13 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U14 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U15 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U16 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U17 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U18 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U19 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U20 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U21 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U22 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U23 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U24 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U25 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U26 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U27 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U28 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U29 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U30 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U31 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U32 (C[59], S[58], X[58], Y[58], Z[58]);
  UBFA_59 U33 (C[60], S[59], X[59], Y[59], Z[59]);
endmodule

module PureCSA_59_30 (C, S, X, Y, Z);
  output [60:31] C;
  output [59:30] S;
  input [59:30] X;
  input [59:30] Y;
  input [59:30] Z;
  UBFA_30 U0 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U1 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U2 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U3 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U4 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U5 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U6 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U7 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U8 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U9 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U10 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U11 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U12 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U13 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U14 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U15 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U16 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U17 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U18 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U19 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U20 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U21 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U22 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U23 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U24 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U25 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U26 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U27 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U28 (C[59], S[58], X[58], Y[58], Z[58]);
  UBFA_59 U29 (C[60], S[59], X[59], Y[59], Z[59]);
endmodule

module PureCSA_62_31 (C, S, X, Y, Z);
  output [63:32] C;
  output [62:31] S;
  input [62:31] X;
  input [62:31] Y;
  input [62:31] Z;
  UBFA_31 U0 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U1 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U2 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U3 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U4 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U5 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U6 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U7 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U8 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U9 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U10 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U11 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U12 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U13 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U14 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U15 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U16 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U17 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U18 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U19 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U20 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U21 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U22 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U23 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U24 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U25 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U26 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U27 (C[59], S[58], X[58], Y[58], Z[58]);
  UBFA_59 U28 (C[60], S[59], X[59], Y[59], Z[59]);
  UBFA_60 U29 (C[61], S[60], X[60], Y[60], Z[60]);
  UBFA_61 U30 (C[62], S[61], X[61], Y[61], Z[61]);
  UBFA_62 U31 (C[63], S[62], X[62], Y[62], Z[62]);
endmodule

module PureCSHA_11_9 (C, S, X, Y);
  output [12:10] C;
  output [11:9] S;
  input [11:9] X;
  input [11:9] Y;
  UBHA_9 U0 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U1 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U2 (C[12], S[11], X[11], Y[11]);
endmodule

module PureCSHA_13_6 (C, S, X, Y);
  output [14:7] C;
  output [13:6] S;
  input [13:6] X;
  input [13:6] Y;
  UBHA_6 U0 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U1 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U2 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U3 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U4 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U5 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U6 (C[13], S[12], X[12], Y[12]);
  UBHA_13 U7 (C[14], S[13], X[13], Y[13]);
endmodule

module PureCSHA_15_13 (C, S, X, Y);
  output [16:14] C;
  output [15:13] S;
  input [15:13] X;
  input [15:13] Y;
  UBHA_13 U0 (C[14], S[13], X[13], Y[13]);
  UBHA_14 U1 (C[15], S[14], X[14], Y[14]);
  UBHA_15 U2 (C[16], S[15], X[15], Y[15]);
endmodule

module PureCSHA_18_7 (C, S, X, Y);
  output [19:8] C;
  output [18:7] S;
  input [18:7] X;
  input [18:7] Y;
  UBHA_7 U0 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U1 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U2 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U3 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U4 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U5 (C[13], S[12], X[12], Y[12]);
  UBHA_13 U6 (C[14], S[13], X[13], Y[13]);
  UBHA_14 U7 (C[15], S[14], X[14], Y[14]);
  UBHA_15 U8 (C[16], S[15], X[15], Y[15]);
  UBHA_16 U9 (C[17], S[16], X[16], Y[16]);
  UBHA_17 U10 (C[18], S[17], X[17], Y[17]);
  UBHA_18 U11 (C[19], S[18], X[18], Y[18]);
endmodule

module PureCSHA_20_18 (C, S, X, Y);
  output [21:19] C;
  output [20:18] S;
  input [20:18] X;
  input [20:18] Y;
  UBHA_18 U0 (C[19], S[18], X[18], Y[18]);
  UBHA_19 U1 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U2 (C[21], S[20], X[20], Y[20]);
endmodule

module PureCSHA_20_19 (C, S, X, Y);
  output [21:20] C;
  output [20:19] S;
  input [20:19] X;
  input [20:19] Y;
  UBHA_19 U0 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U1 (C[21], S[20], X[20], Y[20]);
endmodule

module PureCSHA_21_20 (C, S, X, Y);
  output [22:21] C;
  output [21:20] S;
  input [21:20] X;
  input [21:20] Y;
  UBHA_20 U0 (C[21], S[20], X[20], Y[20]);
  UBHA_21 U1 (C[22], S[21], X[21], Y[21]);
endmodule

module PureCSHA_25_8 (C, S, X, Y);
  output [26:9] C;
  output [25:8] S;
  input [25:8] X;
  input [25:8] Y;
  UBHA_8 U0 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U1 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U2 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U3 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U4 (C[13], S[12], X[12], Y[12]);
  UBHA_13 U5 (C[14], S[13], X[13], Y[13]);
  UBHA_14 U6 (C[15], S[14], X[14], Y[14]);
  UBHA_15 U7 (C[16], S[15], X[15], Y[15]);
  UBHA_16 U8 (C[17], S[16], X[16], Y[16]);
  UBHA_17 U9 (C[18], S[17], X[17], Y[17]);
  UBHA_18 U10 (C[19], S[18], X[18], Y[18]);
  UBHA_19 U11 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U12 (C[21], S[20], X[20], Y[20]);
  UBHA_21 U13 (C[22], S[21], X[21], Y[21]);
  UBHA_22 U14 (C[23], S[22], X[22], Y[22]);
  UBHA_23 U15 (C[24], S[23], X[23], Y[23]);
  UBHA_24 U16 (C[25], S[24], X[24], Y[24]);
  UBHA_25 U17 (C[26], S[25], X[25], Y[25]);
endmodule

module PureCSHA_28_25 (C, S, X, Y);
  output [29:26] C;
  output [28:25] S;
  input [28:25] X;
  input [28:25] Y;
  UBHA_25 U0 (C[26], S[25], X[25], Y[25]);
  UBHA_26 U1 (C[27], S[26], X[26], Y[26]);
  UBHA_27 U2 (C[28], S[27], X[27], Y[27]);
  UBHA_28 U3 (C[29], S[28], X[28], Y[28]);
endmodule

module PureCSHA_28_27 (C, S, X, Y);
  output [29:28] C;
  output [28:27] S;
  input [28:27] X;
  input [28:27] Y;
  UBHA_27 U0 (C[28], S[27], X[27], Y[27]);
  UBHA_28 U1 (C[29], S[28], X[28], Y[28]);
endmodule

module PureCSHA_29_28 (C, S, X, Y);
  output [30:29] C;
  output [29:28] S;
  input [29:28] X;
  input [29:28] Y;
  UBHA_28 U0 (C[29], S[28], X[28], Y[28]);
  UBHA_29 U1 (C[30], S[29], X[29], Y[29]);
endmodule

module PureCSHA_30_28 (C, S, X, Y);
  output [31:29] C;
  output [30:28] S;
  input [30:28] X;
  input [30:28] Y;
  UBHA_28 U0 (C[29], S[28], X[28], Y[28]);
  UBHA_29 U1 (C[30], S[29], X[29], Y[29]);
  UBHA_30 U2 (C[31], S[30], X[30], Y[30]);
endmodule

module PureCSHA_36_35 (C, S, X, Y);
  output [37:36] C;
  output [36:35] S;
  input [36:35] X;
  input [36:35] Y;
  UBHA_35 U0 (C[36], S[35], X[35], Y[35]);
  UBHA_36 U1 (C[37], S[36], X[36], Y[36]);
endmodule

module PureCSHA_39_37 (C, S, X, Y);
  output [40:38] C;
  output [39:37] S;
  input [39:37] X;
  input [39:37] Y;
  UBHA_37 U0 (C[38], S[37], X[37], Y[37]);
  UBHA_38 U1 (C[39], S[38], X[38], Y[38]);
  UBHA_39 U2 (C[40], S[39], X[39], Y[39]);
endmodule

module PureCSHA_39_38 (C, S, X, Y);
  output [40:39] C;
  output [39:38] S;
  input [39:38] X;
  input [39:38] Y;
  UBHA_38 U0 (C[39], S[38], X[38], Y[38]);
  UBHA_39 U1 (C[40], S[39], X[39], Y[39]);
endmodule

module PureCSHA_43_41 (C, S, X, Y);
  output [44:42] C;
  output [43:41] S;
  input [43:41] X;
  input [43:41] Y;
  UBHA_41 U0 (C[42], S[41], X[41], Y[41]);
  UBHA_42 U1 (C[43], S[42], X[42], Y[42]);
  UBHA_43 U2 (C[44], S[43], X[43], Y[43]);
endmodule

module PureCSHA_47_45 (C, S, X, Y);
  output [48:46] C;
  output [47:45] S;
  input [47:45] X;
  input [47:45] Y;
  UBHA_45 U0 (C[46], S[45], X[45], Y[45]);
  UBHA_46 U1 (C[47], S[46], X[46], Y[46]);
  UBHA_47 U2 (C[48], S[47], X[47], Y[47]);
endmodule

module PureCSHA_49_45 (C, S, X, Y);
  output [50:46] C;
  output [49:45] S;
  input [49:45] X;
  input [49:45] Y;
  UBHA_45 U0 (C[46], S[45], X[45], Y[45]);
  UBHA_46 U1 (C[47], S[46], X[46], Y[46]);
  UBHA_47 U2 (C[48], S[47], X[47], Y[47]);
  UBHA_48 U3 (C[49], S[48], X[48], Y[48]);
  UBHA_49 U4 (C[50], S[49], X[49], Y[49]);
endmodule

module PureCSHA_4_3 (C, S, X, Y);
  output [5:4] C;
  output [4:3] S;
  input [4:3] X;
  input [4:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
endmodule

module PureCSHA_52_50 (C, S, X, Y);
  output [53:51] C;
  output [52:50] S;
  input [52:50] X;
  input [52:50] Y;
  UBHA_50 U0 (C[51], S[50], X[50], Y[50]);
  UBHA_51 U1 (C[52], S[51], X[51], Y[51]);
  UBHA_52 U2 (C[53], S[52], X[52], Y[52]);
endmodule

module PureCSHA_54_49 (C, S, X, Y);
  output [55:50] C;
  output [54:49] S;
  input [54:49] X;
  input [54:49] Y;
  UBHA_49 U0 (C[50], S[49], X[49], Y[49]);
  UBHA_50 U1 (C[51], S[50], X[50], Y[50]);
  UBHA_51 U2 (C[52], S[51], X[51], Y[51]);
  UBHA_52 U3 (C[53], S[52], X[52], Y[52]);
  UBHA_53 U4 (C[54], S[53], X[53], Y[53]);
  UBHA_54 U5 (C[55], S[54], X[54], Y[54]);
endmodule

module PureCSHA_58_51 (C, S, X, Y);
  output [59:52] C;
  output [58:51] S;
  input [58:51] X;
  input [58:51] Y;
  UBHA_51 U0 (C[52], S[51], X[51], Y[51]);
  UBHA_52 U1 (C[53], S[52], X[52], Y[52]);
  UBHA_53 U2 (C[54], S[53], X[53], Y[53]);
  UBHA_54 U3 (C[55], S[54], X[54], Y[54]);
  UBHA_55 U4 (C[56], S[55], X[55], Y[55]);
  UBHA_56 U5 (C[57], S[56], X[56], Y[56]);
  UBHA_57 U6 (C[58], S[57], X[57], Y[57]);
  UBHA_58 U7 (C[59], S[58], X[58], Y[58]);
endmodule

module PureCSHA_61_57 (C, S, X, Y);
  output [62:58] C;
  output [61:57] S;
  input [61:57] X;
  input [61:57] Y;
  UBHA_57 U0 (C[58], S[57], X[57], Y[57]);
  UBHA_58 U1 (C[59], S[58], X[58], Y[58]);
  UBHA_59 U2 (C[60], S[59], X[59], Y[59]);
  UBHA_60 U3 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U4 (C[62], S[61], X[61], Y[61]);
endmodule

module PureCSHA_61_59 (C, S, X, Y);
  output [62:60] C;
  output [61:59] S;
  input [61:59] X;
  input [61:59] Y;
  UBHA_59 U0 (C[60], S[59], X[59], Y[59]);
  UBHA_60 U1 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U2 (C[62], S[61], X[61], Y[61]);
endmodule

module PureCSHA_62_56 (C, S, X, Y);
  output [63:57] C;
  output [62:56] S;
  input [62:56] X;
  input [62:56] Y;
  UBHA_56 U0 (C[57], S[56], X[56], Y[56]);
  UBHA_57 U1 (C[58], S[57], X[57], Y[57]);
  UBHA_58 U2 (C[59], S[58], X[58], Y[58]);
  UBHA_59 U3 (C[60], S[59], X[59], Y[59]);
  UBHA_60 U4 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U5 (C[62], S[61], X[61], Y[61]);
  UBHA_62 U6 (C[63], S[62], X[62], Y[62]);
endmodule

module PureCSHA_63_60 (C, S, X, Y);
  output [64:61] C;
  output [63:60] S;
  input [63:60] X;
  input [63:60] Y;
  UBHA_60 U0 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U1 (C[62], S[61], X[61], Y[61]);
  UBHA_62 U2 (C[63], S[62], X[62], Y[62]);
  UBHA_63 U3 (C[64], S[63], X[63], Y[63]);
endmodule

module PureCSHA_6_4 (C, S, X, Y);
  output [7:5] C;
  output [6:4] S;
  input [6:4] X;
  input [6:4] Y;
  UBHA_4 U0 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U1 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U2 (C[7], S[6], X[6], Y[6]);
endmodule

module PureCSHA_7_6 (C, S, X, Y);
  output [8:7] C;
  output [7:6] S;
  input [7:6] X;
  input [7:6] Y;
  UBHA_6 U0 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U1 (C[8], S[7], X[7], Y[7]);
endmodule

module PureCSHA_9_5 (C, S, X, Y);
  output [10:6] C;
  output [9:5] S;
  input [9:5] X;
  input [9:5] Y;
  UBHA_5 U0 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U1 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U2 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U3 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U4 (C[10], S[9], X[9], Y[9]);
endmodule

module TCNVPPG_31_0_31 (O, IN1, IN2);
  output [62:31] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire [61:31] NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UN1BPPG_0_31 U1 (NEG[31], IN1P[0], IN2);
  UN1BPPG_1_31 U2 (NEG[32], IN1P[1], IN2);
  UN1BPPG_2_31 U3 (NEG[33], IN1P[2], IN2);
  UN1BPPG_3_31 U4 (NEG[34], IN1P[3], IN2);
  UN1BPPG_4_31 U5 (NEG[35], IN1P[4], IN2);
  UN1BPPG_5_31 U6 (NEG[36], IN1P[5], IN2);
  UN1BPPG_6_31 U7 (NEG[37], IN1P[6], IN2);
  UN1BPPG_7_31 U8 (NEG[38], IN1P[7], IN2);
  UN1BPPG_8_31 U9 (NEG[39], IN1P[8], IN2);
  UN1BPPG_9_31 U10 (NEG[40], IN1P[9], IN2);
  UN1BPPG_10_31 U11 (NEG[41], IN1P[10], IN2);
  UN1BPPG_11_31 U12 (NEG[42], IN1P[11], IN2);
  UN1BPPG_12_31 U13 (NEG[43], IN1P[12], IN2);
  UN1BPPG_13_31 U14 (NEG[44], IN1P[13], IN2);
  UN1BPPG_14_31 U15 (NEG[45], IN1P[14], IN2);
  UN1BPPG_15_31 U16 (NEG[46], IN1P[15], IN2);
  UN1BPPG_16_31 U17 (NEG[47], IN1P[16], IN2);
  UN1BPPG_17_31 U18 (NEG[48], IN1P[17], IN2);
  UN1BPPG_18_31 U19 (NEG[49], IN1P[18], IN2);
  UN1BPPG_19_31 U20 (NEG[50], IN1P[19], IN2);
  UN1BPPG_20_31 U21 (NEG[51], IN1P[20], IN2);
  UN1BPPG_21_31 U22 (NEG[52], IN1P[21], IN2);
  UN1BPPG_22_31 U23 (NEG[53], IN1P[22], IN2);
  UN1BPPG_23_31 U24 (NEG[54], IN1P[23], IN2);
  UN1BPPG_24_31 U25 (NEG[55], IN1P[24], IN2);
  UN1BPPG_25_31 U26 (NEG[56], IN1P[25], IN2);
  UN1BPPG_26_31 U27 (NEG[57], IN1P[26], IN2);
  UN1BPPG_27_31 U28 (NEG[58], IN1P[27], IN2);
  UN1BPPG_28_31 U29 (NEG[59], IN1P[28], IN2);
  UN1BPPG_29_31 U30 (NEG[60], IN1P[29], IN2);
  UN1BPPG_30_31 U31 (NEG[61], IN1P[30], IN2);
  NUB1BPPG_31_31 U32 (O[62], IN1N, IN2);
  NUBUBCON_61_31 U33 (O[61:31], NEG);
endmodule

module TCPPG_31_0_31_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, IN1, IN2);
  output [32:0] PP0;
  output [32:1] PP1;
  output [41:10] PP10;
  output [42:11] PP11;
  output [43:12] PP12;
  output [44:13] PP13;
  output [45:14] PP14;
  output [46:15] PP15;
  output [47:16] PP16;
  output [48:17] PP17;
  output [49:18] PP18;
  output [50:19] PP19;
  output [33:2] PP2;
  output [51:20] PP20;
  output [52:21] PP21;
  output [53:22] PP22;
  output [54:23] PP23;
  output [55:24] PP24;
  output [56:25] PP25;
  output [57:26] PP26;
  output [58:27] PP27;
  output [59:28] PP28;
  output [60:29] PP29;
  output [34:3] PP3;
  output [61:30] PP30;
  output [62:31] PP31;
  output [35:4] PP4;
  output [36:5] PP5;
  output [37:6] PP6;
  output [38:7] PP7;
  output [39:8] PP8;
  output [40:9] PP9;
  input [31:0] IN1;
  input [31:0] IN2;
  wire BIAS;
  wire [30:0] IN2R;
  wire IN2T;
  wire [31:0] W;
  TCDECON_31_0 U0 (IN2T, IN2R, IN2);
  TCUVPPG_31_0_0 U1 (W, IN1, IN2R[0]);
  TCUVPPG_31_0_1 U2 (PP1, IN1, IN2R[1]);
  TCUVPPG_31_0_2 U3 (PP2, IN1, IN2R[2]);
  TCUVPPG_31_0_3 U4 (PP3, IN1, IN2R[3]);
  TCUVPPG_31_0_4 U5 (PP4, IN1, IN2R[4]);
  TCUVPPG_31_0_5 U6 (PP5, IN1, IN2R[5]);
  TCUVPPG_31_0_6 U7 (PP6, IN1, IN2R[6]);
  TCUVPPG_31_0_7 U8 (PP7, IN1, IN2R[7]);
  TCUVPPG_31_0_8 U9 (PP8, IN1, IN2R[8]);
  TCUVPPG_31_0_9 U10 (PP9, IN1, IN2R[9]);
  TCUVPPG_31_0_10 U11 (PP10, IN1, IN2R[10]);
  TCUVPPG_31_0_11 U12 (PP11, IN1, IN2R[11]);
  TCUVPPG_31_0_12 U13 (PP12, IN1, IN2R[12]);
  TCUVPPG_31_0_13 U14 (PP13, IN1, IN2R[13]);
  TCUVPPG_31_0_14 U15 (PP14, IN1, IN2R[14]);
  TCUVPPG_31_0_15 U16 (PP15, IN1, IN2R[15]);
  TCUVPPG_31_0_16 U17 (PP16, IN1, IN2R[16]);
  TCUVPPG_31_0_17 U18 (PP17, IN1, IN2R[17]);
  TCUVPPG_31_0_18 U19 (PP18, IN1, IN2R[18]);
  TCUVPPG_31_0_19 U20 (PP19, IN1, IN2R[19]);
  TCUVPPG_31_0_20 U21 (PP20, IN1, IN2R[20]);
  TCUVPPG_31_0_21 U22 (PP21, IN1, IN2R[21]);
  TCUVPPG_31_0_22 U23 (PP22, IN1, IN2R[22]);
  TCUVPPG_31_0_23 U24 (PP23, IN1, IN2R[23]);
  TCUVPPG_31_0_24 U25 (PP24, IN1, IN2R[24]);
  TCUVPPG_31_0_25 U26 (PP25, IN1, IN2R[25]);
  TCUVPPG_31_0_26 U27 (PP26, IN1, IN2R[26]);
  TCUVPPG_31_0_27 U28 (PP27, IN1, IN2R[27]);
  TCUVPPG_31_0_28 U29 (PP28, IN1, IN2R[28]);
  TCUVPPG_31_0_29 U30 (PP29, IN1, IN2R[29]);
  TCUVPPG_31_0_30 U31 (PP30, IN1, IN2R[30]);
  TCNVPPG_31_0_31 U32 (PP31, IN1, IN2T);
  UBOne_32 U33 (BIAS);
  UBCMBIN_32_32_31_000 U34 (PP0, BIAS, W);
endmodule

module TCUVPPG_31_0_0 (O, IN1, IN2);
  output [31:0] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_0 U1 (O[0], IN1P[0], IN2);
  UB1BPPG_1_0 U2 (O[1], IN1P[1], IN2);
  UB1BPPG_2_0 U3 (O[2], IN1P[2], IN2);
  UB1BPPG_3_0 U4 (O[3], IN1P[3], IN2);
  UB1BPPG_4_0 U5 (O[4], IN1P[4], IN2);
  UB1BPPG_5_0 U6 (O[5], IN1P[5], IN2);
  UB1BPPG_6_0 U7 (O[6], IN1P[6], IN2);
  UB1BPPG_7_0 U8 (O[7], IN1P[7], IN2);
  UB1BPPG_8_0 U9 (O[8], IN1P[8], IN2);
  UB1BPPG_9_0 U10 (O[9], IN1P[9], IN2);
  UB1BPPG_10_0 U11 (O[10], IN1P[10], IN2);
  UB1BPPG_11_0 U12 (O[11], IN1P[11], IN2);
  UB1BPPG_12_0 U13 (O[12], IN1P[12], IN2);
  UB1BPPG_13_0 U14 (O[13], IN1P[13], IN2);
  UB1BPPG_14_0 U15 (O[14], IN1P[14], IN2);
  UB1BPPG_15_0 U16 (O[15], IN1P[15], IN2);
  UB1BPPG_16_0 U17 (O[16], IN1P[16], IN2);
  UB1BPPG_17_0 U18 (O[17], IN1P[17], IN2);
  UB1BPPG_18_0 U19 (O[18], IN1P[18], IN2);
  UB1BPPG_19_0 U20 (O[19], IN1P[19], IN2);
  UB1BPPG_20_0 U21 (O[20], IN1P[20], IN2);
  UB1BPPG_21_0 U22 (O[21], IN1P[21], IN2);
  UB1BPPG_22_0 U23 (O[22], IN1P[22], IN2);
  UB1BPPG_23_0 U24 (O[23], IN1P[23], IN2);
  UB1BPPG_24_0 U25 (O[24], IN1P[24], IN2);
  UB1BPPG_25_0 U26 (O[25], IN1P[25], IN2);
  UB1BPPG_26_0 U27 (O[26], IN1P[26], IN2);
  UB1BPPG_27_0 U28 (O[27], IN1P[27], IN2);
  UB1BPPG_28_0 U29 (O[28], IN1P[28], IN2);
  UB1BPPG_29_0 U30 (O[29], IN1P[29], IN2);
  UB1BPPG_30_0 U31 (O[30], IN1P[30], IN2);
  NU1BPPG_31_0 U32 (NEG, IN1N, IN2);
  NUBUB1CON_31 U33 (O[31], NEG);
endmodule

module TCUVPPG_31_0_1 (O, IN1, IN2);
  output [32:1] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_1 U1 (O[1], IN1P[0], IN2);
  UB1BPPG_1_1 U2 (O[2], IN1P[1], IN2);
  UB1BPPG_2_1 U3 (O[3], IN1P[2], IN2);
  UB1BPPG_3_1 U4 (O[4], IN1P[3], IN2);
  UB1BPPG_4_1 U5 (O[5], IN1P[4], IN2);
  UB1BPPG_5_1 U6 (O[6], IN1P[5], IN2);
  UB1BPPG_6_1 U7 (O[7], IN1P[6], IN2);
  UB1BPPG_7_1 U8 (O[8], IN1P[7], IN2);
  UB1BPPG_8_1 U9 (O[9], IN1P[8], IN2);
  UB1BPPG_9_1 U10 (O[10], IN1P[9], IN2);
  UB1BPPG_10_1 U11 (O[11], IN1P[10], IN2);
  UB1BPPG_11_1 U12 (O[12], IN1P[11], IN2);
  UB1BPPG_12_1 U13 (O[13], IN1P[12], IN2);
  UB1BPPG_13_1 U14 (O[14], IN1P[13], IN2);
  UB1BPPG_14_1 U15 (O[15], IN1P[14], IN2);
  UB1BPPG_15_1 U16 (O[16], IN1P[15], IN2);
  UB1BPPG_16_1 U17 (O[17], IN1P[16], IN2);
  UB1BPPG_17_1 U18 (O[18], IN1P[17], IN2);
  UB1BPPG_18_1 U19 (O[19], IN1P[18], IN2);
  UB1BPPG_19_1 U20 (O[20], IN1P[19], IN2);
  UB1BPPG_20_1 U21 (O[21], IN1P[20], IN2);
  UB1BPPG_21_1 U22 (O[22], IN1P[21], IN2);
  UB1BPPG_22_1 U23 (O[23], IN1P[22], IN2);
  UB1BPPG_23_1 U24 (O[24], IN1P[23], IN2);
  UB1BPPG_24_1 U25 (O[25], IN1P[24], IN2);
  UB1BPPG_25_1 U26 (O[26], IN1P[25], IN2);
  UB1BPPG_26_1 U27 (O[27], IN1P[26], IN2);
  UB1BPPG_27_1 U28 (O[28], IN1P[27], IN2);
  UB1BPPG_28_1 U29 (O[29], IN1P[28], IN2);
  UB1BPPG_29_1 U30 (O[30], IN1P[29], IN2);
  UB1BPPG_30_1 U31 (O[31], IN1P[30], IN2);
  NU1BPPG_31_1 U32 (NEG, IN1N, IN2);
  NUBUB1CON_32 U33 (O[32], NEG);
endmodule

module TCUVPPG_31_0_10 (O, IN1, IN2);
  output [41:10] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_10 U1 (O[10], IN1P[0], IN2);
  UB1BPPG_1_10 U2 (O[11], IN1P[1], IN2);
  UB1BPPG_2_10 U3 (O[12], IN1P[2], IN2);
  UB1BPPG_3_10 U4 (O[13], IN1P[3], IN2);
  UB1BPPG_4_10 U5 (O[14], IN1P[4], IN2);
  UB1BPPG_5_10 U6 (O[15], IN1P[5], IN2);
  UB1BPPG_6_10 U7 (O[16], IN1P[6], IN2);
  UB1BPPG_7_10 U8 (O[17], IN1P[7], IN2);
  UB1BPPG_8_10 U9 (O[18], IN1P[8], IN2);
  UB1BPPG_9_10 U10 (O[19], IN1P[9], IN2);
  UB1BPPG_10_10 U11 (O[20], IN1P[10], IN2);
  UB1BPPG_11_10 U12 (O[21], IN1P[11], IN2);
  UB1BPPG_12_10 U13 (O[22], IN1P[12], IN2);
  UB1BPPG_13_10 U14 (O[23], IN1P[13], IN2);
  UB1BPPG_14_10 U15 (O[24], IN1P[14], IN2);
  UB1BPPG_15_10 U16 (O[25], IN1P[15], IN2);
  UB1BPPG_16_10 U17 (O[26], IN1P[16], IN2);
  UB1BPPG_17_10 U18 (O[27], IN1P[17], IN2);
  UB1BPPG_18_10 U19 (O[28], IN1P[18], IN2);
  UB1BPPG_19_10 U20 (O[29], IN1P[19], IN2);
  UB1BPPG_20_10 U21 (O[30], IN1P[20], IN2);
  UB1BPPG_21_10 U22 (O[31], IN1P[21], IN2);
  UB1BPPG_22_10 U23 (O[32], IN1P[22], IN2);
  UB1BPPG_23_10 U24 (O[33], IN1P[23], IN2);
  UB1BPPG_24_10 U25 (O[34], IN1P[24], IN2);
  UB1BPPG_25_10 U26 (O[35], IN1P[25], IN2);
  UB1BPPG_26_10 U27 (O[36], IN1P[26], IN2);
  UB1BPPG_27_10 U28 (O[37], IN1P[27], IN2);
  UB1BPPG_28_10 U29 (O[38], IN1P[28], IN2);
  UB1BPPG_29_10 U30 (O[39], IN1P[29], IN2);
  UB1BPPG_30_10 U31 (O[40], IN1P[30], IN2);
  NU1BPPG_31_10 U32 (NEG, IN1N, IN2);
  NUBUB1CON_41 U33 (O[41], NEG);
endmodule

module TCUVPPG_31_0_11 (O, IN1, IN2);
  output [42:11] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_11 U1 (O[11], IN1P[0], IN2);
  UB1BPPG_1_11 U2 (O[12], IN1P[1], IN2);
  UB1BPPG_2_11 U3 (O[13], IN1P[2], IN2);
  UB1BPPG_3_11 U4 (O[14], IN1P[3], IN2);
  UB1BPPG_4_11 U5 (O[15], IN1P[4], IN2);
  UB1BPPG_5_11 U6 (O[16], IN1P[5], IN2);
  UB1BPPG_6_11 U7 (O[17], IN1P[6], IN2);
  UB1BPPG_7_11 U8 (O[18], IN1P[7], IN2);
  UB1BPPG_8_11 U9 (O[19], IN1P[8], IN2);
  UB1BPPG_9_11 U10 (O[20], IN1P[9], IN2);
  UB1BPPG_10_11 U11 (O[21], IN1P[10], IN2);
  UB1BPPG_11_11 U12 (O[22], IN1P[11], IN2);
  UB1BPPG_12_11 U13 (O[23], IN1P[12], IN2);
  UB1BPPG_13_11 U14 (O[24], IN1P[13], IN2);
  UB1BPPG_14_11 U15 (O[25], IN1P[14], IN2);
  UB1BPPG_15_11 U16 (O[26], IN1P[15], IN2);
  UB1BPPG_16_11 U17 (O[27], IN1P[16], IN2);
  UB1BPPG_17_11 U18 (O[28], IN1P[17], IN2);
  UB1BPPG_18_11 U19 (O[29], IN1P[18], IN2);
  UB1BPPG_19_11 U20 (O[30], IN1P[19], IN2);
  UB1BPPG_20_11 U21 (O[31], IN1P[20], IN2);
  UB1BPPG_21_11 U22 (O[32], IN1P[21], IN2);
  UB1BPPG_22_11 U23 (O[33], IN1P[22], IN2);
  UB1BPPG_23_11 U24 (O[34], IN1P[23], IN2);
  UB1BPPG_24_11 U25 (O[35], IN1P[24], IN2);
  UB1BPPG_25_11 U26 (O[36], IN1P[25], IN2);
  UB1BPPG_26_11 U27 (O[37], IN1P[26], IN2);
  UB1BPPG_27_11 U28 (O[38], IN1P[27], IN2);
  UB1BPPG_28_11 U29 (O[39], IN1P[28], IN2);
  UB1BPPG_29_11 U30 (O[40], IN1P[29], IN2);
  UB1BPPG_30_11 U31 (O[41], IN1P[30], IN2);
  NU1BPPG_31_11 U32 (NEG, IN1N, IN2);
  NUBUB1CON_42 U33 (O[42], NEG);
endmodule

module TCUVPPG_31_0_12 (O, IN1, IN2);
  output [43:12] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_12 U1 (O[12], IN1P[0], IN2);
  UB1BPPG_1_12 U2 (O[13], IN1P[1], IN2);
  UB1BPPG_2_12 U3 (O[14], IN1P[2], IN2);
  UB1BPPG_3_12 U4 (O[15], IN1P[3], IN2);
  UB1BPPG_4_12 U5 (O[16], IN1P[4], IN2);
  UB1BPPG_5_12 U6 (O[17], IN1P[5], IN2);
  UB1BPPG_6_12 U7 (O[18], IN1P[6], IN2);
  UB1BPPG_7_12 U8 (O[19], IN1P[7], IN2);
  UB1BPPG_8_12 U9 (O[20], IN1P[8], IN2);
  UB1BPPG_9_12 U10 (O[21], IN1P[9], IN2);
  UB1BPPG_10_12 U11 (O[22], IN1P[10], IN2);
  UB1BPPG_11_12 U12 (O[23], IN1P[11], IN2);
  UB1BPPG_12_12 U13 (O[24], IN1P[12], IN2);
  UB1BPPG_13_12 U14 (O[25], IN1P[13], IN2);
  UB1BPPG_14_12 U15 (O[26], IN1P[14], IN2);
  UB1BPPG_15_12 U16 (O[27], IN1P[15], IN2);
  UB1BPPG_16_12 U17 (O[28], IN1P[16], IN2);
  UB1BPPG_17_12 U18 (O[29], IN1P[17], IN2);
  UB1BPPG_18_12 U19 (O[30], IN1P[18], IN2);
  UB1BPPG_19_12 U20 (O[31], IN1P[19], IN2);
  UB1BPPG_20_12 U21 (O[32], IN1P[20], IN2);
  UB1BPPG_21_12 U22 (O[33], IN1P[21], IN2);
  UB1BPPG_22_12 U23 (O[34], IN1P[22], IN2);
  UB1BPPG_23_12 U24 (O[35], IN1P[23], IN2);
  UB1BPPG_24_12 U25 (O[36], IN1P[24], IN2);
  UB1BPPG_25_12 U26 (O[37], IN1P[25], IN2);
  UB1BPPG_26_12 U27 (O[38], IN1P[26], IN2);
  UB1BPPG_27_12 U28 (O[39], IN1P[27], IN2);
  UB1BPPG_28_12 U29 (O[40], IN1P[28], IN2);
  UB1BPPG_29_12 U30 (O[41], IN1P[29], IN2);
  UB1BPPG_30_12 U31 (O[42], IN1P[30], IN2);
  NU1BPPG_31_12 U32 (NEG, IN1N, IN2);
  NUBUB1CON_43 U33 (O[43], NEG);
endmodule

module TCUVPPG_31_0_13 (O, IN1, IN2);
  output [44:13] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_13 U1 (O[13], IN1P[0], IN2);
  UB1BPPG_1_13 U2 (O[14], IN1P[1], IN2);
  UB1BPPG_2_13 U3 (O[15], IN1P[2], IN2);
  UB1BPPG_3_13 U4 (O[16], IN1P[3], IN2);
  UB1BPPG_4_13 U5 (O[17], IN1P[4], IN2);
  UB1BPPG_5_13 U6 (O[18], IN1P[5], IN2);
  UB1BPPG_6_13 U7 (O[19], IN1P[6], IN2);
  UB1BPPG_7_13 U8 (O[20], IN1P[7], IN2);
  UB1BPPG_8_13 U9 (O[21], IN1P[8], IN2);
  UB1BPPG_9_13 U10 (O[22], IN1P[9], IN2);
  UB1BPPG_10_13 U11 (O[23], IN1P[10], IN2);
  UB1BPPG_11_13 U12 (O[24], IN1P[11], IN2);
  UB1BPPG_12_13 U13 (O[25], IN1P[12], IN2);
  UB1BPPG_13_13 U14 (O[26], IN1P[13], IN2);
  UB1BPPG_14_13 U15 (O[27], IN1P[14], IN2);
  UB1BPPG_15_13 U16 (O[28], IN1P[15], IN2);
  UB1BPPG_16_13 U17 (O[29], IN1P[16], IN2);
  UB1BPPG_17_13 U18 (O[30], IN1P[17], IN2);
  UB1BPPG_18_13 U19 (O[31], IN1P[18], IN2);
  UB1BPPG_19_13 U20 (O[32], IN1P[19], IN2);
  UB1BPPG_20_13 U21 (O[33], IN1P[20], IN2);
  UB1BPPG_21_13 U22 (O[34], IN1P[21], IN2);
  UB1BPPG_22_13 U23 (O[35], IN1P[22], IN2);
  UB1BPPG_23_13 U24 (O[36], IN1P[23], IN2);
  UB1BPPG_24_13 U25 (O[37], IN1P[24], IN2);
  UB1BPPG_25_13 U26 (O[38], IN1P[25], IN2);
  UB1BPPG_26_13 U27 (O[39], IN1P[26], IN2);
  UB1BPPG_27_13 U28 (O[40], IN1P[27], IN2);
  UB1BPPG_28_13 U29 (O[41], IN1P[28], IN2);
  UB1BPPG_29_13 U30 (O[42], IN1P[29], IN2);
  UB1BPPG_30_13 U31 (O[43], IN1P[30], IN2);
  NU1BPPG_31_13 U32 (NEG, IN1N, IN2);
  NUBUB1CON_44 U33 (O[44], NEG);
endmodule

module TCUVPPG_31_0_14 (O, IN1, IN2);
  output [45:14] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_14 U1 (O[14], IN1P[0], IN2);
  UB1BPPG_1_14 U2 (O[15], IN1P[1], IN2);
  UB1BPPG_2_14 U3 (O[16], IN1P[2], IN2);
  UB1BPPG_3_14 U4 (O[17], IN1P[3], IN2);
  UB1BPPG_4_14 U5 (O[18], IN1P[4], IN2);
  UB1BPPG_5_14 U6 (O[19], IN1P[5], IN2);
  UB1BPPG_6_14 U7 (O[20], IN1P[6], IN2);
  UB1BPPG_7_14 U8 (O[21], IN1P[7], IN2);
  UB1BPPG_8_14 U9 (O[22], IN1P[8], IN2);
  UB1BPPG_9_14 U10 (O[23], IN1P[9], IN2);
  UB1BPPG_10_14 U11 (O[24], IN1P[10], IN2);
  UB1BPPG_11_14 U12 (O[25], IN1P[11], IN2);
  UB1BPPG_12_14 U13 (O[26], IN1P[12], IN2);
  UB1BPPG_13_14 U14 (O[27], IN1P[13], IN2);
  UB1BPPG_14_14 U15 (O[28], IN1P[14], IN2);
  UB1BPPG_15_14 U16 (O[29], IN1P[15], IN2);
  UB1BPPG_16_14 U17 (O[30], IN1P[16], IN2);
  UB1BPPG_17_14 U18 (O[31], IN1P[17], IN2);
  UB1BPPG_18_14 U19 (O[32], IN1P[18], IN2);
  UB1BPPG_19_14 U20 (O[33], IN1P[19], IN2);
  UB1BPPG_20_14 U21 (O[34], IN1P[20], IN2);
  UB1BPPG_21_14 U22 (O[35], IN1P[21], IN2);
  UB1BPPG_22_14 U23 (O[36], IN1P[22], IN2);
  UB1BPPG_23_14 U24 (O[37], IN1P[23], IN2);
  UB1BPPG_24_14 U25 (O[38], IN1P[24], IN2);
  UB1BPPG_25_14 U26 (O[39], IN1P[25], IN2);
  UB1BPPG_26_14 U27 (O[40], IN1P[26], IN2);
  UB1BPPG_27_14 U28 (O[41], IN1P[27], IN2);
  UB1BPPG_28_14 U29 (O[42], IN1P[28], IN2);
  UB1BPPG_29_14 U30 (O[43], IN1P[29], IN2);
  UB1BPPG_30_14 U31 (O[44], IN1P[30], IN2);
  NU1BPPG_31_14 U32 (NEG, IN1N, IN2);
  NUBUB1CON_45 U33 (O[45], NEG);
endmodule

module TCUVPPG_31_0_15 (O, IN1, IN2);
  output [46:15] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_15 U1 (O[15], IN1P[0], IN2);
  UB1BPPG_1_15 U2 (O[16], IN1P[1], IN2);
  UB1BPPG_2_15 U3 (O[17], IN1P[2], IN2);
  UB1BPPG_3_15 U4 (O[18], IN1P[3], IN2);
  UB1BPPG_4_15 U5 (O[19], IN1P[4], IN2);
  UB1BPPG_5_15 U6 (O[20], IN1P[5], IN2);
  UB1BPPG_6_15 U7 (O[21], IN1P[6], IN2);
  UB1BPPG_7_15 U8 (O[22], IN1P[7], IN2);
  UB1BPPG_8_15 U9 (O[23], IN1P[8], IN2);
  UB1BPPG_9_15 U10 (O[24], IN1P[9], IN2);
  UB1BPPG_10_15 U11 (O[25], IN1P[10], IN2);
  UB1BPPG_11_15 U12 (O[26], IN1P[11], IN2);
  UB1BPPG_12_15 U13 (O[27], IN1P[12], IN2);
  UB1BPPG_13_15 U14 (O[28], IN1P[13], IN2);
  UB1BPPG_14_15 U15 (O[29], IN1P[14], IN2);
  UB1BPPG_15_15 U16 (O[30], IN1P[15], IN2);
  UB1BPPG_16_15 U17 (O[31], IN1P[16], IN2);
  UB1BPPG_17_15 U18 (O[32], IN1P[17], IN2);
  UB1BPPG_18_15 U19 (O[33], IN1P[18], IN2);
  UB1BPPG_19_15 U20 (O[34], IN1P[19], IN2);
  UB1BPPG_20_15 U21 (O[35], IN1P[20], IN2);
  UB1BPPG_21_15 U22 (O[36], IN1P[21], IN2);
  UB1BPPG_22_15 U23 (O[37], IN1P[22], IN2);
  UB1BPPG_23_15 U24 (O[38], IN1P[23], IN2);
  UB1BPPG_24_15 U25 (O[39], IN1P[24], IN2);
  UB1BPPG_25_15 U26 (O[40], IN1P[25], IN2);
  UB1BPPG_26_15 U27 (O[41], IN1P[26], IN2);
  UB1BPPG_27_15 U28 (O[42], IN1P[27], IN2);
  UB1BPPG_28_15 U29 (O[43], IN1P[28], IN2);
  UB1BPPG_29_15 U30 (O[44], IN1P[29], IN2);
  UB1BPPG_30_15 U31 (O[45], IN1P[30], IN2);
  NU1BPPG_31_15 U32 (NEG, IN1N, IN2);
  NUBUB1CON_46 U33 (O[46], NEG);
endmodule

module TCUVPPG_31_0_16 (O, IN1, IN2);
  output [47:16] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_16 U1 (O[16], IN1P[0], IN2);
  UB1BPPG_1_16 U2 (O[17], IN1P[1], IN2);
  UB1BPPG_2_16 U3 (O[18], IN1P[2], IN2);
  UB1BPPG_3_16 U4 (O[19], IN1P[3], IN2);
  UB1BPPG_4_16 U5 (O[20], IN1P[4], IN2);
  UB1BPPG_5_16 U6 (O[21], IN1P[5], IN2);
  UB1BPPG_6_16 U7 (O[22], IN1P[6], IN2);
  UB1BPPG_7_16 U8 (O[23], IN1P[7], IN2);
  UB1BPPG_8_16 U9 (O[24], IN1P[8], IN2);
  UB1BPPG_9_16 U10 (O[25], IN1P[9], IN2);
  UB1BPPG_10_16 U11 (O[26], IN1P[10], IN2);
  UB1BPPG_11_16 U12 (O[27], IN1P[11], IN2);
  UB1BPPG_12_16 U13 (O[28], IN1P[12], IN2);
  UB1BPPG_13_16 U14 (O[29], IN1P[13], IN2);
  UB1BPPG_14_16 U15 (O[30], IN1P[14], IN2);
  UB1BPPG_15_16 U16 (O[31], IN1P[15], IN2);
  UB1BPPG_16_16 U17 (O[32], IN1P[16], IN2);
  UB1BPPG_17_16 U18 (O[33], IN1P[17], IN2);
  UB1BPPG_18_16 U19 (O[34], IN1P[18], IN2);
  UB1BPPG_19_16 U20 (O[35], IN1P[19], IN2);
  UB1BPPG_20_16 U21 (O[36], IN1P[20], IN2);
  UB1BPPG_21_16 U22 (O[37], IN1P[21], IN2);
  UB1BPPG_22_16 U23 (O[38], IN1P[22], IN2);
  UB1BPPG_23_16 U24 (O[39], IN1P[23], IN2);
  UB1BPPG_24_16 U25 (O[40], IN1P[24], IN2);
  UB1BPPG_25_16 U26 (O[41], IN1P[25], IN2);
  UB1BPPG_26_16 U27 (O[42], IN1P[26], IN2);
  UB1BPPG_27_16 U28 (O[43], IN1P[27], IN2);
  UB1BPPG_28_16 U29 (O[44], IN1P[28], IN2);
  UB1BPPG_29_16 U30 (O[45], IN1P[29], IN2);
  UB1BPPG_30_16 U31 (O[46], IN1P[30], IN2);
  NU1BPPG_31_16 U32 (NEG, IN1N, IN2);
  NUBUB1CON_47 U33 (O[47], NEG);
endmodule

module TCUVPPG_31_0_17 (O, IN1, IN2);
  output [48:17] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_17 U1 (O[17], IN1P[0], IN2);
  UB1BPPG_1_17 U2 (O[18], IN1P[1], IN2);
  UB1BPPG_2_17 U3 (O[19], IN1P[2], IN2);
  UB1BPPG_3_17 U4 (O[20], IN1P[3], IN2);
  UB1BPPG_4_17 U5 (O[21], IN1P[4], IN2);
  UB1BPPG_5_17 U6 (O[22], IN1P[5], IN2);
  UB1BPPG_6_17 U7 (O[23], IN1P[6], IN2);
  UB1BPPG_7_17 U8 (O[24], IN1P[7], IN2);
  UB1BPPG_8_17 U9 (O[25], IN1P[8], IN2);
  UB1BPPG_9_17 U10 (O[26], IN1P[9], IN2);
  UB1BPPG_10_17 U11 (O[27], IN1P[10], IN2);
  UB1BPPG_11_17 U12 (O[28], IN1P[11], IN2);
  UB1BPPG_12_17 U13 (O[29], IN1P[12], IN2);
  UB1BPPG_13_17 U14 (O[30], IN1P[13], IN2);
  UB1BPPG_14_17 U15 (O[31], IN1P[14], IN2);
  UB1BPPG_15_17 U16 (O[32], IN1P[15], IN2);
  UB1BPPG_16_17 U17 (O[33], IN1P[16], IN2);
  UB1BPPG_17_17 U18 (O[34], IN1P[17], IN2);
  UB1BPPG_18_17 U19 (O[35], IN1P[18], IN2);
  UB1BPPG_19_17 U20 (O[36], IN1P[19], IN2);
  UB1BPPG_20_17 U21 (O[37], IN1P[20], IN2);
  UB1BPPG_21_17 U22 (O[38], IN1P[21], IN2);
  UB1BPPG_22_17 U23 (O[39], IN1P[22], IN2);
  UB1BPPG_23_17 U24 (O[40], IN1P[23], IN2);
  UB1BPPG_24_17 U25 (O[41], IN1P[24], IN2);
  UB1BPPG_25_17 U26 (O[42], IN1P[25], IN2);
  UB1BPPG_26_17 U27 (O[43], IN1P[26], IN2);
  UB1BPPG_27_17 U28 (O[44], IN1P[27], IN2);
  UB1BPPG_28_17 U29 (O[45], IN1P[28], IN2);
  UB1BPPG_29_17 U30 (O[46], IN1P[29], IN2);
  UB1BPPG_30_17 U31 (O[47], IN1P[30], IN2);
  NU1BPPG_31_17 U32 (NEG, IN1N, IN2);
  NUBUB1CON_48 U33 (O[48], NEG);
endmodule

module TCUVPPG_31_0_18 (O, IN1, IN2);
  output [49:18] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_18 U1 (O[18], IN1P[0], IN2);
  UB1BPPG_1_18 U2 (O[19], IN1P[1], IN2);
  UB1BPPG_2_18 U3 (O[20], IN1P[2], IN2);
  UB1BPPG_3_18 U4 (O[21], IN1P[3], IN2);
  UB1BPPG_4_18 U5 (O[22], IN1P[4], IN2);
  UB1BPPG_5_18 U6 (O[23], IN1P[5], IN2);
  UB1BPPG_6_18 U7 (O[24], IN1P[6], IN2);
  UB1BPPG_7_18 U8 (O[25], IN1P[7], IN2);
  UB1BPPG_8_18 U9 (O[26], IN1P[8], IN2);
  UB1BPPG_9_18 U10 (O[27], IN1P[9], IN2);
  UB1BPPG_10_18 U11 (O[28], IN1P[10], IN2);
  UB1BPPG_11_18 U12 (O[29], IN1P[11], IN2);
  UB1BPPG_12_18 U13 (O[30], IN1P[12], IN2);
  UB1BPPG_13_18 U14 (O[31], IN1P[13], IN2);
  UB1BPPG_14_18 U15 (O[32], IN1P[14], IN2);
  UB1BPPG_15_18 U16 (O[33], IN1P[15], IN2);
  UB1BPPG_16_18 U17 (O[34], IN1P[16], IN2);
  UB1BPPG_17_18 U18 (O[35], IN1P[17], IN2);
  UB1BPPG_18_18 U19 (O[36], IN1P[18], IN2);
  UB1BPPG_19_18 U20 (O[37], IN1P[19], IN2);
  UB1BPPG_20_18 U21 (O[38], IN1P[20], IN2);
  UB1BPPG_21_18 U22 (O[39], IN1P[21], IN2);
  UB1BPPG_22_18 U23 (O[40], IN1P[22], IN2);
  UB1BPPG_23_18 U24 (O[41], IN1P[23], IN2);
  UB1BPPG_24_18 U25 (O[42], IN1P[24], IN2);
  UB1BPPG_25_18 U26 (O[43], IN1P[25], IN2);
  UB1BPPG_26_18 U27 (O[44], IN1P[26], IN2);
  UB1BPPG_27_18 U28 (O[45], IN1P[27], IN2);
  UB1BPPG_28_18 U29 (O[46], IN1P[28], IN2);
  UB1BPPG_29_18 U30 (O[47], IN1P[29], IN2);
  UB1BPPG_30_18 U31 (O[48], IN1P[30], IN2);
  NU1BPPG_31_18 U32 (NEG, IN1N, IN2);
  NUBUB1CON_49 U33 (O[49], NEG);
endmodule

module TCUVPPG_31_0_19 (O, IN1, IN2);
  output [50:19] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_19 U1 (O[19], IN1P[0], IN2);
  UB1BPPG_1_19 U2 (O[20], IN1P[1], IN2);
  UB1BPPG_2_19 U3 (O[21], IN1P[2], IN2);
  UB1BPPG_3_19 U4 (O[22], IN1P[3], IN2);
  UB1BPPG_4_19 U5 (O[23], IN1P[4], IN2);
  UB1BPPG_5_19 U6 (O[24], IN1P[5], IN2);
  UB1BPPG_6_19 U7 (O[25], IN1P[6], IN2);
  UB1BPPG_7_19 U8 (O[26], IN1P[7], IN2);
  UB1BPPG_8_19 U9 (O[27], IN1P[8], IN2);
  UB1BPPG_9_19 U10 (O[28], IN1P[9], IN2);
  UB1BPPG_10_19 U11 (O[29], IN1P[10], IN2);
  UB1BPPG_11_19 U12 (O[30], IN1P[11], IN2);
  UB1BPPG_12_19 U13 (O[31], IN1P[12], IN2);
  UB1BPPG_13_19 U14 (O[32], IN1P[13], IN2);
  UB1BPPG_14_19 U15 (O[33], IN1P[14], IN2);
  UB1BPPG_15_19 U16 (O[34], IN1P[15], IN2);
  UB1BPPG_16_19 U17 (O[35], IN1P[16], IN2);
  UB1BPPG_17_19 U18 (O[36], IN1P[17], IN2);
  UB1BPPG_18_19 U19 (O[37], IN1P[18], IN2);
  UB1BPPG_19_19 U20 (O[38], IN1P[19], IN2);
  UB1BPPG_20_19 U21 (O[39], IN1P[20], IN2);
  UB1BPPG_21_19 U22 (O[40], IN1P[21], IN2);
  UB1BPPG_22_19 U23 (O[41], IN1P[22], IN2);
  UB1BPPG_23_19 U24 (O[42], IN1P[23], IN2);
  UB1BPPG_24_19 U25 (O[43], IN1P[24], IN2);
  UB1BPPG_25_19 U26 (O[44], IN1P[25], IN2);
  UB1BPPG_26_19 U27 (O[45], IN1P[26], IN2);
  UB1BPPG_27_19 U28 (O[46], IN1P[27], IN2);
  UB1BPPG_28_19 U29 (O[47], IN1P[28], IN2);
  UB1BPPG_29_19 U30 (O[48], IN1P[29], IN2);
  UB1BPPG_30_19 U31 (O[49], IN1P[30], IN2);
  NU1BPPG_31_19 U32 (NEG, IN1N, IN2);
  NUBUB1CON_50 U33 (O[50], NEG);
endmodule

module TCUVPPG_31_0_2 (O, IN1, IN2);
  output [33:2] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_2 U1 (O[2], IN1P[0], IN2);
  UB1BPPG_1_2 U2 (O[3], IN1P[1], IN2);
  UB1BPPG_2_2 U3 (O[4], IN1P[2], IN2);
  UB1BPPG_3_2 U4 (O[5], IN1P[3], IN2);
  UB1BPPG_4_2 U5 (O[6], IN1P[4], IN2);
  UB1BPPG_5_2 U6 (O[7], IN1P[5], IN2);
  UB1BPPG_6_2 U7 (O[8], IN1P[6], IN2);
  UB1BPPG_7_2 U8 (O[9], IN1P[7], IN2);
  UB1BPPG_8_2 U9 (O[10], IN1P[8], IN2);
  UB1BPPG_9_2 U10 (O[11], IN1P[9], IN2);
  UB1BPPG_10_2 U11 (O[12], IN1P[10], IN2);
  UB1BPPG_11_2 U12 (O[13], IN1P[11], IN2);
  UB1BPPG_12_2 U13 (O[14], IN1P[12], IN2);
  UB1BPPG_13_2 U14 (O[15], IN1P[13], IN2);
  UB1BPPG_14_2 U15 (O[16], IN1P[14], IN2);
  UB1BPPG_15_2 U16 (O[17], IN1P[15], IN2);
  UB1BPPG_16_2 U17 (O[18], IN1P[16], IN2);
  UB1BPPG_17_2 U18 (O[19], IN1P[17], IN2);
  UB1BPPG_18_2 U19 (O[20], IN1P[18], IN2);
  UB1BPPG_19_2 U20 (O[21], IN1P[19], IN2);
  UB1BPPG_20_2 U21 (O[22], IN1P[20], IN2);
  UB1BPPG_21_2 U22 (O[23], IN1P[21], IN2);
  UB1BPPG_22_2 U23 (O[24], IN1P[22], IN2);
  UB1BPPG_23_2 U24 (O[25], IN1P[23], IN2);
  UB1BPPG_24_2 U25 (O[26], IN1P[24], IN2);
  UB1BPPG_25_2 U26 (O[27], IN1P[25], IN2);
  UB1BPPG_26_2 U27 (O[28], IN1P[26], IN2);
  UB1BPPG_27_2 U28 (O[29], IN1P[27], IN2);
  UB1BPPG_28_2 U29 (O[30], IN1P[28], IN2);
  UB1BPPG_29_2 U30 (O[31], IN1P[29], IN2);
  UB1BPPG_30_2 U31 (O[32], IN1P[30], IN2);
  NU1BPPG_31_2 U32 (NEG, IN1N, IN2);
  NUBUB1CON_33 U33 (O[33], NEG);
endmodule

module TCUVPPG_31_0_20 (O, IN1, IN2);
  output [51:20] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_20 U1 (O[20], IN1P[0], IN2);
  UB1BPPG_1_20 U2 (O[21], IN1P[1], IN2);
  UB1BPPG_2_20 U3 (O[22], IN1P[2], IN2);
  UB1BPPG_3_20 U4 (O[23], IN1P[3], IN2);
  UB1BPPG_4_20 U5 (O[24], IN1P[4], IN2);
  UB1BPPG_5_20 U6 (O[25], IN1P[5], IN2);
  UB1BPPG_6_20 U7 (O[26], IN1P[6], IN2);
  UB1BPPG_7_20 U8 (O[27], IN1P[7], IN2);
  UB1BPPG_8_20 U9 (O[28], IN1P[8], IN2);
  UB1BPPG_9_20 U10 (O[29], IN1P[9], IN2);
  UB1BPPG_10_20 U11 (O[30], IN1P[10], IN2);
  UB1BPPG_11_20 U12 (O[31], IN1P[11], IN2);
  UB1BPPG_12_20 U13 (O[32], IN1P[12], IN2);
  UB1BPPG_13_20 U14 (O[33], IN1P[13], IN2);
  UB1BPPG_14_20 U15 (O[34], IN1P[14], IN2);
  UB1BPPG_15_20 U16 (O[35], IN1P[15], IN2);
  UB1BPPG_16_20 U17 (O[36], IN1P[16], IN2);
  UB1BPPG_17_20 U18 (O[37], IN1P[17], IN2);
  UB1BPPG_18_20 U19 (O[38], IN1P[18], IN2);
  UB1BPPG_19_20 U20 (O[39], IN1P[19], IN2);
  UB1BPPG_20_20 U21 (O[40], IN1P[20], IN2);
  UB1BPPG_21_20 U22 (O[41], IN1P[21], IN2);
  UB1BPPG_22_20 U23 (O[42], IN1P[22], IN2);
  UB1BPPG_23_20 U24 (O[43], IN1P[23], IN2);
  UB1BPPG_24_20 U25 (O[44], IN1P[24], IN2);
  UB1BPPG_25_20 U26 (O[45], IN1P[25], IN2);
  UB1BPPG_26_20 U27 (O[46], IN1P[26], IN2);
  UB1BPPG_27_20 U28 (O[47], IN1P[27], IN2);
  UB1BPPG_28_20 U29 (O[48], IN1P[28], IN2);
  UB1BPPG_29_20 U30 (O[49], IN1P[29], IN2);
  UB1BPPG_30_20 U31 (O[50], IN1P[30], IN2);
  NU1BPPG_31_20 U32 (NEG, IN1N, IN2);
  NUBUB1CON_51 U33 (O[51], NEG);
endmodule

module TCUVPPG_31_0_21 (O, IN1, IN2);
  output [52:21] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_21 U1 (O[21], IN1P[0], IN2);
  UB1BPPG_1_21 U2 (O[22], IN1P[1], IN2);
  UB1BPPG_2_21 U3 (O[23], IN1P[2], IN2);
  UB1BPPG_3_21 U4 (O[24], IN1P[3], IN2);
  UB1BPPG_4_21 U5 (O[25], IN1P[4], IN2);
  UB1BPPG_5_21 U6 (O[26], IN1P[5], IN2);
  UB1BPPG_6_21 U7 (O[27], IN1P[6], IN2);
  UB1BPPG_7_21 U8 (O[28], IN1P[7], IN2);
  UB1BPPG_8_21 U9 (O[29], IN1P[8], IN2);
  UB1BPPG_9_21 U10 (O[30], IN1P[9], IN2);
  UB1BPPG_10_21 U11 (O[31], IN1P[10], IN2);
  UB1BPPG_11_21 U12 (O[32], IN1P[11], IN2);
  UB1BPPG_12_21 U13 (O[33], IN1P[12], IN2);
  UB1BPPG_13_21 U14 (O[34], IN1P[13], IN2);
  UB1BPPG_14_21 U15 (O[35], IN1P[14], IN2);
  UB1BPPG_15_21 U16 (O[36], IN1P[15], IN2);
  UB1BPPG_16_21 U17 (O[37], IN1P[16], IN2);
  UB1BPPG_17_21 U18 (O[38], IN1P[17], IN2);
  UB1BPPG_18_21 U19 (O[39], IN1P[18], IN2);
  UB1BPPG_19_21 U20 (O[40], IN1P[19], IN2);
  UB1BPPG_20_21 U21 (O[41], IN1P[20], IN2);
  UB1BPPG_21_21 U22 (O[42], IN1P[21], IN2);
  UB1BPPG_22_21 U23 (O[43], IN1P[22], IN2);
  UB1BPPG_23_21 U24 (O[44], IN1P[23], IN2);
  UB1BPPG_24_21 U25 (O[45], IN1P[24], IN2);
  UB1BPPG_25_21 U26 (O[46], IN1P[25], IN2);
  UB1BPPG_26_21 U27 (O[47], IN1P[26], IN2);
  UB1BPPG_27_21 U28 (O[48], IN1P[27], IN2);
  UB1BPPG_28_21 U29 (O[49], IN1P[28], IN2);
  UB1BPPG_29_21 U30 (O[50], IN1P[29], IN2);
  UB1BPPG_30_21 U31 (O[51], IN1P[30], IN2);
  NU1BPPG_31_21 U32 (NEG, IN1N, IN2);
  NUBUB1CON_52 U33 (O[52], NEG);
endmodule

module TCUVPPG_31_0_22 (O, IN1, IN2);
  output [53:22] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_22 U1 (O[22], IN1P[0], IN2);
  UB1BPPG_1_22 U2 (O[23], IN1P[1], IN2);
  UB1BPPG_2_22 U3 (O[24], IN1P[2], IN2);
  UB1BPPG_3_22 U4 (O[25], IN1P[3], IN2);
  UB1BPPG_4_22 U5 (O[26], IN1P[4], IN2);
  UB1BPPG_5_22 U6 (O[27], IN1P[5], IN2);
  UB1BPPG_6_22 U7 (O[28], IN1P[6], IN2);
  UB1BPPG_7_22 U8 (O[29], IN1P[7], IN2);
  UB1BPPG_8_22 U9 (O[30], IN1P[8], IN2);
  UB1BPPG_9_22 U10 (O[31], IN1P[9], IN2);
  UB1BPPG_10_22 U11 (O[32], IN1P[10], IN2);
  UB1BPPG_11_22 U12 (O[33], IN1P[11], IN2);
  UB1BPPG_12_22 U13 (O[34], IN1P[12], IN2);
  UB1BPPG_13_22 U14 (O[35], IN1P[13], IN2);
  UB1BPPG_14_22 U15 (O[36], IN1P[14], IN2);
  UB1BPPG_15_22 U16 (O[37], IN1P[15], IN2);
  UB1BPPG_16_22 U17 (O[38], IN1P[16], IN2);
  UB1BPPG_17_22 U18 (O[39], IN1P[17], IN2);
  UB1BPPG_18_22 U19 (O[40], IN1P[18], IN2);
  UB1BPPG_19_22 U20 (O[41], IN1P[19], IN2);
  UB1BPPG_20_22 U21 (O[42], IN1P[20], IN2);
  UB1BPPG_21_22 U22 (O[43], IN1P[21], IN2);
  UB1BPPG_22_22 U23 (O[44], IN1P[22], IN2);
  UB1BPPG_23_22 U24 (O[45], IN1P[23], IN2);
  UB1BPPG_24_22 U25 (O[46], IN1P[24], IN2);
  UB1BPPG_25_22 U26 (O[47], IN1P[25], IN2);
  UB1BPPG_26_22 U27 (O[48], IN1P[26], IN2);
  UB1BPPG_27_22 U28 (O[49], IN1P[27], IN2);
  UB1BPPG_28_22 U29 (O[50], IN1P[28], IN2);
  UB1BPPG_29_22 U30 (O[51], IN1P[29], IN2);
  UB1BPPG_30_22 U31 (O[52], IN1P[30], IN2);
  NU1BPPG_31_22 U32 (NEG, IN1N, IN2);
  NUBUB1CON_53 U33 (O[53], NEG);
endmodule

module TCUVPPG_31_0_23 (O, IN1, IN2);
  output [54:23] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_23 U1 (O[23], IN1P[0], IN2);
  UB1BPPG_1_23 U2 (O[24], IN1P[1], IN2);
  UB1BPPG_2_23 U3 (O[25], IN1P[2], IN2);
  UB1BPPG_3_23 U4 (O[26], IN1P[3], IN2);
  UB1BPPG_4_23 U5 (O[27], IN1P[4], IN2);
  UB1BPPG_5_23 U6 (O[28], IN1P[5], IN2);
  UB1BPPG_6_23 U7 (O[29], IN1P[6], IN2);
  UB1BPPG_7_23 U8 (O[30], IN1P[7], IN2);
  UB1BPPG_8_23 U9 (O[31], IN1P[8], IN2);
  UB1BPPG_9_23 U10 (O[32], IN1P[9], IN2);
  UB1BPPG_10_23 U11 (O[33], IN1P[10], IN2);
  UB1BPPG_11_23 U12 (O[34], IN1P[11], IN2);
  UB1BPPG_12_23 U13 (O[35], IN1P[12], IN2);
  UB1BPPG_13_23 U14 (O[36], IN1P[13], IN2);
  UB1BPPG_14_23 U15 (O[37], IN1P[14], IN2);
  UB1BPPG_15_23 U16 (O[38], IN1P[15], IN2);
  UB1BPPG_16_23 U17 (O[39], IN1P[16], IN2);
  UB1BPPG_17_23 U18 (O[40], IN1P[17], IN2);
  UB1BPPG_18_23 U19 (O[41], IN1P[18], IN2);
  UB1BPPG_19_23 U20 (O[42], IN1P[19], IN2);
  UB1BPPG_20_23 U21 (O[43], IN1P[20], IN2);
  UB1BPPG_21_23 U22 (O[44], IN1P[21], IN2);
  UB1BPPG_22_23 U23 (O[45], IN1P[22], IN2);
  UB1BPPG_23_23 U24 (O[46], IN1P[23], IN2);
  UB1BPPG_24_23 U25 (O[47], IN1P[24], IN2);
  UB1BPPG_25_23 U26 (O[48], IN1P[25], IN2);
  UB1BPPG_26_23 U27 (O[49], IN1P[26], IN2);
  UB1BPPG_27_23 U28 (O[50], IN1P[27], IN2);
  UB1BPPG_28_23 U29 (O[51], IN1P[28], IN2);
  UB1BPPG_29_23 U30 (O[52], IN1P[29], IN2);
  UB1BPPG_30_23 U31 (O[53], IN1P[30], IN2);
  NU1BPPG_31_23 U32 (NEG, IN1N, IN2);
  NUBUB1CON_54 U33 (O[54], NEG);
endmodule

module TCUVPPG_31_0_24 (O, IN1, IN2);
  output [55:24] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_24 U1 (O[24], IN1P[0], IN2);
  UB1BPPG_1_24 U2 (O[25], IN1P[1], IN2);
  UB1BPPG_2_24 U3 (O[26], IN1P[2], IN2);
  UB1BPPG_3_24 U4 (O[27], IN1P[3], IN2);
  UB1BPPG_4_24 U5 (O[28], IN1P[4], IN2);
  UB1BPPG_5_24 U6 (O[29], IN1P[5], IN2);
  UB1BPPG_6_24 U7 (O[30], IN1P[6], IN2);
  UB1BPPG_7_24 U8 (O[31], IN1P[7], IN2);
  UB1BPPG_8_24 U9 (O[32], IN1P[8], IN2);
  UB1BPPG_9_24 U10 (O[33], IN1P[9], IN2);
  UB1BPPG_10_24 U11 (O[34], IN1P[10], IN2);
  UB1BPPG_11_24 U12 (O[35], IN1P[11], IN2);
  UB1BPPG_12_24 U13 (O[36], IN1P[12], IN2);
  UB1BPPG_13_24 U14 (O[37], IN1P[13], IN2);
  UB1BPPG_14_24 U15 (O[38], IN1P[14], IN2);
  UB1BPPG_15_24 U16 (O[39], IN1P[15], IN2);
  UB1BPPG_16_24 U17 (O[40], IN1P[16], IN2);
  UB1BPPG_17_24 U18 (O[41], IN1P[17], IN2);
  UB1BPPG_18_24 U19 (O[42], IN1P[18], IN2);
  UB1BPPG_19_24 U20 (O[43], IN1P[19], IN2);
  UB1BPPG_20_24 U21 (O[44], IN1P[20], IN2);
  UB1BPPG_21_24 U22 (O[45], IN1P[21], IN2);
  UB1BPPG_22_24 U23 (O[46], IN1P[22], IN2);
  UB1BPPG_23_24 U24 (O[47], IN1P[23], IN2);
  UB1BPPG_24_24 U25 (O[48], IN1P[24], IN2);
  UB1BPPG_25_24 U26 (O[49], IN1P[25], IN2);
  UB1BPPG_26_24 U27 (O[50], IN1P[26], IN2);
  UB1BPPG_27_24 U28 (O[51], IN1P[27], IN2);
  UB1BPPG_28_24 U29 (O[52], IN1P[28], IN2);
  UB1BPPG_29_24 U30 (O[53], IN1P[29], IN2);
  UB1BPPG_30_24 U31 (O[54], IN1P[30], IN2);
  NU1BPPG_31_24 U32 (NEG, IN1N, IN2);
  NUBUB1CON_55 U33 (O[55], NEG);
endmodule

module TCUVPPG_31_0_25 (O, IN1, IN2);
  output [56:25] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_25 U1 (O[25], IN1P[0], IN2);
  UB1BPPG_1_25 U2 (O[26], IN1P[1], IN2);
  UB1BPPG_2_25 U3 (O[27], IN1P[2], IN2);
  UB1BPPG_3_25 U4 (O[28], IN1P[3], IN2);
  UB1BPPG_4_25 U5 (O[29], IN1P[4], IN2);
  UB1BPPG_5_25 U6 (O[30], IN1P[5], IN2);
  UB1BPPG_6_25 U7 (O[31], IN1P[6], IN2);
  UB1BPPG_7_25 U8 (O[32], IN1P[7], IN2);
  UB1BPPG_8_25 U9 (O[33], IN1P[8], IN2);
  UB1BPPG_9_25 U10 (O[34], IN1P[9], IN2);
  UB1BPPG_10_25 U11 (O[35], IN1P[10], IN2);
  UB1BPPG_11_25 U12 (O[36], IN1P[11], IN2);
  UB1BPPG_12_25 U13 (O[37], IN1P[12], IN2);
  UB1BPPG_13_25 U14 (O[38], IN1P[13], IN2);
  UB1BPPG_14_25 U15 (O[39], IN1P[14], IN2);
  UB1BPPG_15_25 U16 (O[40], IN1P[15], IN2);
  UB1BPPG_16_25 U17 (O[41], IN1P[16], IN2);
  UB1BPPG_17_25 U18 (O[42], IN1P[17], IN2);
  UB1BPPG_18_25 U19 (O[43], IN1P[18], IN2);
  UB1BPPG_19_25 U20 (O[44], IN1P[19], IN2);
  UB1BPPG_20_25 U21 (O[45], IN1P[20], IN2);
  UB1BPPG_21_25 U22 (O[46], IN1P[21], IN2);
  UB1BPPG_22_25 U23 (O[47], IN1P[22], IN2);
  UB1BPPG_23_25 U24 (O[48], IN1P[23], IN2);
  UB1BPPG_24_25 U25 (O[49], IN1P[24], IN2);
  UB1BPPG_25_25 U26 (O[50], IN1P[25], IN2);
  UB1BPPG_26_25 U27 (O[51], IN1P[26], IN2);
  UB1BPPG_27_25 U28 (O[52], IN1P[27], IN2);
  UB1BPPG_28_25 U29 (O[53], IN1P[28], IN2);
  UB1BPPG_29_25 U30 (O[54], IN1P[29], IN2);
  UB1BPPG_30_25 U31 (O[55], IN1P[30], IN2);
  NU1BPPG_31_25 U32 (NEG, IN1N, IN2);
  NUBUB1CON_56 U33 (O[56], NEG);
endmodule

module TCUVPPG_31_0_26 (O, IN1, IN2);
  output [57:26] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_26 U1 (O[26], IN1P[0], IN2);
  UB1BPPG_1_26 U2 (O[27], IN1P[1], IN2);
  UB1BPPG_2_26 U3 (O[28], IN1P[2], IN2);
  UB1BPPG_3_26 U4 (O[29], IN1P[3], IN2);
  UB1BPPG_4_26 U5 (O[30], IN1P[4], IN2);
  UB1BPPG_5_26 U6 (O[31], IN1P[5], IN2);
  UB1BPPG_6_26 U7 (O[32], IN1P[6], IN2);
  UB1BPPG_7_26 U8 (O[33], IN1P[7], IN2);
  UB1BPPG_8_26 U9 (O[34], IN1P[8], IN2);
  UB1BPPG_9_26 U10 (O[35], IN1P[9], IN2);
  UB1BPPG_10_26 U11 (O[36], IN1P[10], IN2);
  UB1BPPG_11_26 U12 (O[37], IN1P[11], IN2);
  UB1BPPG_12_26 U13 (O[38], IN1P[12], IN2);
  UB1BPPG_13_26 U14 (O[39], IN1P[13], IN2);
  UB1BPPG_14_26 U15 (O[40], IN1P[14], IN2);
  UB1BPPG_15_26 U16 (O[41], IN1P[15], IN2);
  UB1BPPG_16_26 U17 (O[42], IN1P[16], IN2);
  UB1BPPG_17_26 U18 (O[43], IN1P[17], IN2);
  UB1BPPG_18_26 U19 (O[44], IN1P[18], IN2);
  UB1BPPG_19_26 U20 (O[45], IN1P[19], IN2);
  UB1BPPG_20_26 U21 (O[46], IN1P[20], IN2);
  UB1BPPG_21_26 U22 (O[47], IN1P[21], IN2);
  UB1BPPG_22_26 U23 (O[48], IN1P[22], IN2);
  UB1BPPG_23_26 U24 (O[49], IN1P[23], IN2);
  UB1BPPG_24_26 U25 (O[50], IN1P[24], IN2);
  UB1BPPG_25_26 U26 (O[51], IN1P[25], IN2);
  UB1BPPG_26_26 U27 (O[52], IN1P[26], IN2);
  UB1BPPG_27_26 U28 (O[53], IN1P[27], IN2);
  UB1BPPG_28_26 U29 (O[54], IN1P[28], IN2);
  UB1BPPG_29_26 U30 (O[55], IN1P[29], IN2);
  UB1BPPG_30_26 U31 (O[56], IN1P[30], IN2);
  NU1BPPG_31_26 U32 (NEG, IN1N, IN2);
  NUBUB1CON_57 U33 (O[57], NEG);
endmodule

module TCUVPPG_31_0_27 (O, IN1, IN2);
  output [58:27] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_27 U1 (O[27], IN1P[0], IN2);
  UB1BPPG_1_27 U2 (O[28], IN1P[1], IN2);
  UB1BPPG_2_27 U3 (O[29], IN1P[2], IN2);
  UB1BPPG_3_27 U4 (O[30], IN1P[3], IN2);
  UB1BPPG_4_27 U5 (O[31], IN1P[4], IN2);
  UB1BPPG_5_27 U6 (O[32], IN1P[5], IN2);
  UB1BPPG_6_27 U7 (O[33], IN1P[6], IN2);
  UB1BPPG_7_27 U8 (O[34], IN1P[7], IN2);
  UB1BPPG_8_27 U9 (O[35], IN1P[8], IN2);
  UB1BPPG_9_27 U10 (O[36], IN1P[9], IN2);
  UB1BPPG_10_27 U11 (O[37], IN1P[10], IN2);
  UB1BPPG_11_27 U12 (O[38], IN1P[11], IN2);
  UB1BPPG_12_27 U13 (O[39], IN1P[12], IN2);
  UB1BPPG_13_27 U14 (O[40], IN1P[13], IN2);
  UB1BPPG_14_27 U15 (O[41], IN1P[14], IN2);
  UB1BPPG_15_27 U16 (O[42], IN1P[15], IN2);
  UB1BPPG_16_27 U17 (O[43], IN1P[16], IN2);
  UB1BPPG_17_27 U18 (O[44], IN1P[17], IN2);
  UB1BPPG_18_27 U19 (O[45], IN1P[18], IN2);
  UB1BPPG_19_27 U20 (O[46], IN1P[19], IN2);
  UB1BPPG_20_27 U21 (O[47], IN1P[20], IN2);
  UB1BPPG_21_27 U22 (O[48], IN1P[21], IN2);
  UB1BPPG_22_27 U23 (O[49], IN1P[22], IN2);
  UB1BPPG_23_27 U24 (O[50], IN1P[23], IN2);
  UB1BPPG_24_27 U25 (O[51], IN1P[24], IN2);
  UB1BPPG_25_27 U26 (O[52], IN1P[25], IN2);
  UB1BPPG_26_27 U27 (O[53], IN1P[26], IN2);
  UB1BPPG_27_27 U28 (O[54], IN1P[27], IN2);
  UB1BPPG_28_27 U29 (O[55], IN1P[28], IN2);
  UB1BPPG_29_27 U30 (O[56], IN1P[29], IN2);
  UB1BPPG_30_27 U31 (O[57], IN1P[30], IN2);
  NU1BPPG_31_27 U32 (NEG, IN1N, IN2);
  NUBUB1CON_58 U33 (O[58], NEG);
endmodule

module TCUVPPG_31_0_28 (O, IN1, IN2);
  output [59:28] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_28 U1 (O[28], IN1P[0], IN2);
  UB1BPPG_1_28 U2 (O[29], IN1P[1], IN2);
  UB1BPPG_2_28 U3 (O[30], IN1P[2], IN2);
  UB1BPPG_3_28 U4 (O[31], IN1P[3], IN2);
  UB1BPPG_4_28 U5 (O[32], IN1P[4], IN2);
  UB1BPPG_5_28 U6 (O[33], IN1P[5], IN2);
  UB1BPPG_6_28 U7 (O[34], IN1P[6], IN2);
  UB1BPPG_7_28 U8 (O[35], IN1P[7], IN2);
  UB1BPPG_8_28 U9 (O[36], IN1P[8], IN2);
  UB1BPPG_9_28 U10 (O[37], IN1P[9], IN2);
  UB1BPPG_10_28 U11 (O[38], IN1P[10], IN2);
  UB1BPPG_11_28 U12 (O[39], IN1P[11], IN2);
  UB1BPPG_12_28 U13 (O[40], IN1P[12], IN2);
  UB1BPPG_13_28 U14 (O[41], IN1P[13], IN2);
  UB1BPPG_14_28 U15 (O[42], IN1P[14], IN2);
  UB1BPPG_15_28 U16 (O[43], IN1P[15], IN2);
  UB1BPPG_16_28 U17 (O[44], IN1P[16], IN2);
  UB1BPPG_17_28 U18 (O[45], IN1P[17], IN2);
  UB1BPPG_18_28 U19 (O[46], IN1P[18], IN2);
  UB1BPPG_19_28 U20 (O[47], IN1P[19], IN2);
  UB1BPPG_20_28 U21 (O[48], IN1P[20], IN2);
  UB1BPPG_21_28 U22 (O[49], IN1P[21], IN2);
  UB1BPPG_22_28 U23 (O[50], IN1P[22], IN2);
  UB1BPPG_23_28 U24 (O[51], IN1P[23], IN2);
  UB1BPPG_24_28 U25 (O[52], IN1P[24], IN2);
  UB1BPPG_25_28 U26 (O[53], IN1P[25], IN2);
  UB1BPPG_26_28 U27 (O[54], IN1P[26], IN2);
  UB1BPPG_27_28 U28 (O[55], IN1P[27], IN2);
  UB1BPPG_28_28 U29 (O[56], IN1P[28], IN2);
  UB1BPPG_29_28 U30 (O[57], IN1P[29], IN2);
  UB1BPPG_30_28 U31 (O[58], IN1P[30], IN2);
  NU1BPPG_31_28 U32 (NEG, IN1N, IN2);
  NUBUB1CON_59 U33 (O[59], NEG);
endmodule

module TCUVPPG_31_0_29 (O, IN1, IN2);
  output [60:29] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_29 U1 (O[29], IN1P[0], IN2);
  UB1BPPG_1_29 U2 (O[30], IN1P[1], IN2);
  UB1BPPG_2_29 U3 (O[31], IN1P[2], IN2);
  UB1BPPG_3_29 U4 (O[32], IN1P[3], IN2);
  UB1BPPG_4_29 U5 (O[33], IN1P[4], IN2);
  UB1BPPG_5_29 U6 (O[34], IN1P[5], IN2);
  UB1BPPG_6_29 U7 (O[35], IN1P[6], IN2);
  UB1BPPG_7_29 U8 (O[36], IN1P[7], IN2);
  UB1BPPG_8_29 U9 (O[37], IN1P[8], IN2);
  UB1BPPG_9_29 U10 (O[38], IN1P[9], IN2);
  UB1BPPG_10_29 U11 (O[39], IN1P[10], IN2);
  UB1BPPG_11_29 U12 (O[40], IN1P[11], IN2);
  UB1BPPG_12_29 U13 (O[41], IN1P[12], IN2);
  UB1BPPG_13_29 U14 (O[42], IN1P[13], IN2);
  UB1BPPG_14_29 U15 (O[43], IN1P[14], IN2);
  UB1BPPG_15_29 U16 (O[44], IN1P[15], IN2);
  UB1BPPG_16_29 U17 (O[45], IN1P[16], IN2);
  UB1BPPG_17_29 U18 (O[46], IN1P[17], IN2);
  UB1BPPG_18_29 U19 (O[47], IN1P[18], IN2);
  UB1BPPG_19_29 U20 (O[48], IN1P[19], IN2);
  UB1BPPG_20_29 U21 (O[49], IN1P[20], IN2);
  UB1BPPG_21_29 U22 (O[50], IN1P[21], IN2);
  UB1BPPG_22_29 U23 (O[51], IN1P[22], IN2);
  UB1BPPG_23_29 U24 (O[52], IN1P[23], IN2);
  UB1BPPG_24_29 U25 (O[53], IN1P[24], IN2);
  UB1BPPG_25_29 U26 (O[54], IN1P[25], IN2);
  UB1BPPG_26_29 U27 (O[55], IN1P[26], IN2);
  UB1BPPG_27_29 U28 (O[56], IN1P[27], IN2);
  UB1BPPG_28_29 U29 (O[57], IN1P[28], IN2);
  UB1BPPG_29_29 U30 (O[58], IN1P[29], IN2);
  UB1BPPG_30_29 U31 (O[59], IN1P[30], IN2);
  NU1BPPG_31_29 U32 (NEG, IN1N, IN2);
  NUBUB1CON_60 U33 (O[60], NEG);
endmodule

module TCUVPPG_31_0_3 (O, IN1, IN2);
  output [34:3] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_3 U1 (O[3], IN1P[0], IN2);
  UB1BPPG_1_3 U2 (O[4], IN1P[1], IN2);
  UB1BPPG_2_3 U3 (O[5], IN1P[2], IN2);
  UB1BPPG_3_3 U4 (O[6], IN1P[3], IN2);
  UB1BPPG_4_3 U5 (O[7], IN1P[4], IN2);
  UB1BPPG_5_3 U6 (O[8], IN1P[5], IN2);
  UB1BPPG_6_3 U7 (O[9], IN1P[6], IN2);
  UB1BPPG_7_3 U8 (O[10], IN1P[7], IN2);
  UB1BPPG_8_3 U9 (O[11], IN1P[8], IN2);
  UB1BPPG_9_3 U10 (O[12], IN1P[9], IN2);
  UB1BPPG_10_3 U11 (O[13], IN1P[10], IN2);
  UB1BPPG_11_3 U12 (O[14], IN1P[11], IN2);
  UB1BPPG_12_3 U13 (O[15], IN1P[12], IN2);
  UB1BPPG_13_3 U14 (O[16], IN1P[13], IN2);
  UB1BPPG_14_3 U15 (O[17], IN1P[14], IN2);
  UB1BPPG_15_3 U16 (O[18], IN1P[15], IN2);
  UB1BPPG_16_3 U17 (O[19], IN1P[16], IN2);
  UB1BPPG_17_3 U18 (O[20], IN1P[17], IN2);
  UB1BPPG_18_3 U19 (O[21], IN1P[18], IN2);
  UB1BPPG_19_3 U20 (O[22], IN1P[19], IN2);
  UB1BPPG_20_3 U21 (O[23], IN1P[20], IN2);
  UB1BPPG_21_3 U22 (O[24], IN1P[21], IN2);
  UB1BPPG_22_3 U23 (O[25], IN1P[22], IN2);
  UB1BPPG_23_3 U24 (O[26], IN1P[23], IN2);
  UB1BPPG_24_3 U25 (O[27], IN1P[24], IN2);
  UB1BPPG_25_3 U26 (O[28], IN1P[25], IN2);
  UB1BPPG_26_3 U27 (O[29], IN1P[26], IN2);
  UB1BPPG_27_3 U28 (O[30], IN1P[27], IN2);
  UB1BPPG_28_3 U29 (O[31], IN1P[28], IN2);
  UB1BPPG_29_3 U30 (O[32], IN1P[29], IN2);
  UB1BPPG_30_3 U31 (O[33], IN1P[30], IN2);
  NU1BPPG_31_3 U32 (NEG, IN1N, IN2);
  NUBUB1CON_34 U33 (O[34], NEG);
endmodule

module TCUVPPG_31_0_30 (O, IN1, IN2);
  output [61:30] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_30 U1 (O[30], IN1P[0], IN2);
  UB1BPPG_1_30 U2 (O[31], IN1P[1], IN2);
  UB1BPPG_2_30 U3 (O[32], IN1P[2], IN2);
  UB1BPPG_3_30 U4 (O[33], IN1P[3], IN2);
  UB1BPPG_4_30 U5 (O[34], IN1P[4], IN2);
  UB1BPPG_5_30 U6 (O[35], IN1P[5], IN2);
  UB1BPPG_6_30 U7 (O[36], IN1P[6], IN2);
  UB1BPPG_7_30 U8 (O[37], IN1P[7], IN2);
  UB1BPPG_8_30 U9 (O[38], IN1P[8], IN2);
  UB1BPPG_9_30 U10 (O[39], IN1P[9], IN2);
  UB1BPPG_10_30 U11 (O[40], IN1P[10], IN2);
  UB1BPPG_11_30 U12 (O[41], IN1P[11], IN2);
  UB1BPPG_12_30 U13 (O[42], IN1P[12], IN2);
  UB1BPPG_13_30 U14 (O[43], IN1P[13], IN2);
  UB1BPPG_14_30 U15 (O[44], IN1P[14], IN2);
  UB1BPPG_15_30 U16 (O[45], IN1P[15], IN2);
  UB1BPPG_16_30 U17 (O[46], IN1P[16], IN2);
  UB1BPPG_17_30 U18 (O[47], IN1P[17], IN2);
  UB1BPPG_18_30 U19 (O[48], IN1P[18], IN2);
  UB1BPPG_19_30 U20 (O[49], IN1P[19], IN2);
  UB1BPPG_20_30 U21 (O[50], IN1P[20], IN2);
  UB1BPPG_21_30 U22 (O[51], IN1P[21], IN2);
  UB1BPPG_22_30 U23 (O[52], IN1P[22], IN2);
  UB1BPPG_23_30 U24 (O[53], IN1P[23], IN2);
  UB1BPPG_24_30 U25 (O[54], IN1P[24], IN2);
  UB1BPPG_25_30 U26 (O[55], IN1P[25], IN2);
  UB1BPPG_26_30 U27 (O[56], IN1P[26], IN2);
  UB1BPPG_27_30 U28 (O[57], IN1P[27], IN2);
  UB1BPPG_28_30 U29 (O[58], IN1P[28], IN2);
  UB1BPPG_29_30 U30 (O[59], IN1P[29], IN2);
  UB1BPPG_30_30 U31 (O[60], IN1P[30], IN2);
  NU1BPPG_31_30 U32 (NEG, IN1N, IN2);
  NUBUB1CON_61 U33 (O[61], NEG);
endmodule

module TCUVPPG_31_0_4 (O, IN1, IN2);
  output [35:4] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_4 U1 (O[4], IN1P[0], IN2);
  UB1BPPG_1_4 U2 (O[5], IN1P[1], IN2);
  UB1BPPG_2_4 U3 (O[6], IN1P[2], IN2);
  UB1BPPG_3_4 U4 (O[7], IN1P[3], IN2);
  UB1BPPG_4_4 U5 (O[8], IN1P[4], IN2);
  UB1BPPG_5_4 U6 (O[9], IN1P[5], IN2);
  UB1BPPG_6_4 U7 (O[10], IN1P[6], IN2);
  UB1BPPG_7_4 U8 (O[11], IN1P[7], IN2);
  UB1BPPG_8_4 U9 (O[12], IN1P[8], IN2);
  UB1BPPG_9_4 U10 (O[13], IN1P[9], IN2);
  UB1BPPG_10_4 U11 (O[14], IN1P[10], IN2);
  UB1BPPG_11_4 U12 (O[15], IN1P[11], IN2);
  UB1BPPG_12_4 U13 (O[16], IN1P[12], IN2);
  UB1BPPG_13_4 U14 (O[17], IN1P[13], IN2);
  UB1BPPG_14_4 U15 (O[18], IN1P[14], IN2);
  UB1BPPG_15_4 U16 (O[19], IN1P[15], IN2);
  UB1BPPG_16_4 U17 (O[20], IN1P[16], IN2);
  UB1BPPG_17_4 U18 (O[21], IN1P[17], IN2);
  UB1BPPG_18_4 U19 (O[22], IN1P[18], IN2);
  UB1BPPG_19_4 U20 (O[23], IN1P[19], IN2);
  UB1BPPG_20_4 U21 (O[24], IN1P[20], IN2);
  UB1BPPG_21_4 U22 (O[25], IN1P[21], IN2);
  UB1BPPG_22_4 U23 (O[26], IN1P[22], IN2);
  UB1BPPG_23_4 U24 (O[27], IN1P[23], IN2);
  UB1BPPG_24_4 U25 (O[28], IN1P[24], IN2);
  UB1BPPG_25_4 U26 (O[29], IN1P[25], IN2);
  UB1BPPG_26_4 U27 (O[30], IN1P[26], IN2);
  UB1BPPG_27_4 U28 (O[31], IN1P[27], IN2);
  UB1BPPG_28_4 U29 (O[32], IN1P[28], IN2);
  UB1BPPG_29_4 U30 (O[33], IN1P[29], IN2);
  UB1BPPG_30_4 U31 (O[34], IN1P[30], IN2);
  NU1BPPG_31_4 U32 (NEG, IN1N, IN2);
  NUBUB1CON_35 U33 (O[35], NEG);
endmodule

module TCUVPPG_31_0_5 (O, IN1, IN2);
  output [36:5] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_5 U1 (O[5], IN1P[0], IN2);
  UB1BPPG_1_5 U2 (O[6], IN1P[1], IN2);
  UB1BPPG_2_5 U3 (O[7], IN1P[2], IN2);
  UB1BPPG_3_5 U4 (O[8], IN1P[3], IN2);
  UB1BPPG_4_5 U5 (O[9], IN1P[4], IN2);
  UB1BPPG_5_5 U6 (O[10], IN1P[5], IN2);
  UB1BPPG_6_5 U7 (O[11], IN1P[6], IN2);
  UB1BPPG_7_5 U8 (O[12], IN1P[7], IN2);
  UB1BPPG_8_5 U9 (O[13], IN1P[8], IN2);
  UB1BPPG_9_5 U10 (O[14], IN1P[9], IN2);
  UB1BPPG_10_5 U11 (O[15], IN1P[10], IN2);
  UB1BPPG_11_5 U12 (O[16], IN1P[11], IN2);
  UB1BPPG_12_5 U13 (O[17], IN1P[12], IN2);
  UB1BPPG_13_5 U14 (O[18], IN1P[13], IN2);
  UB1BPPG_14_5 U15 (O[19], IN1P[14], IN2);
  UB1BPPG_15_5 U16 (O[20], IN1P[15], IN2);
  UB1BPPG_16_5 U17 (O[21], IN1P[16], IN2);
  UB1BPPG_17_5 U18 (O[22], IN1P[17], IN2);
  UB1BPPG_18_5 U19 (O[23], IN1P[18], IN2);
  UB1BPPG_19_5 U20 (O[24], IN1P[19], IN2);
  UB1BPPG_20_5 U21 (O[25], IN1P[20], IN2);
  UB1BPPG_21_5 U22 (O[26], IN1P[21], IN2);
  UB1BPPG_22_5 U23 (O[27], IN1P[22], IN2);
  UB1BPPG_23_5 U24 (O[28], IN1P[23], IN2);
  UB1BPPG_24_5 U25 (O[29], IN1P[24], IN2);
  UB1BPPG_25_5 U26 (O[30], IN1P[25], IN2);
  UB1BPPG_26_5 U27 (O[31], IN1P[26], IN2);
  UB1BPPG_27_5 U28 (O[32], IN1P[27], IN2);
  UB1BPPG_28_5 U29 (O[33], IN1P[28], IN2);
  UB1BPPG_29_5 U30 (O[34], IN1P[29], IN2);
  UB1BPPG_30_5 U31 (O[35], IN1P[30], IN2);
  NU1BPPG_31_5 U32 (NEG, IN1N, IN2);
  NUBUB1CON_36 U33 (O[36], NEG);
endmodule

module TCUVPPG_31_0_6 (O, IN1, IN2);
  output [37:6] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_6 U1 (O[6], IN1P[0], IN2);
  UB1BPPG_1_6 U2 (O[7], IN1P[1], IN2);
  UB1BPPG_2_6 U3 (O[8], IN1P[2], IN2);
  UB1BPPG_3_6 U4 (O[9], IN1P[3], IN2);
  UB1BPPG_4_6 U5 (O[10], IN1P[4], IN2);
  UB1BPPG_5_6 U6 (O[11], IN1P[5], IN2);
  UB1BPPG_6_6 U7 (O[12], IN1P[6], IN2);
  UB1BPPG_7_6 U8 (O[13], IN1P[7], IN2);
  UB1BPPG_8_6 U9 (O[14], IN1P[8], IN2);
  UB1BPPG_9_6 U10 (O[15], IN1P[9], IN2);
  UB1BPPG_10_6 U11 (O[16], IN1P[10], IN2);
  UB1BPPG_11_6 U12 (O[17], IN1P[11], IN2);
  UB1BPPG_12_6 U13 (O[18], IN1P[12], IN2);
  UB1BPPG_13_6 U14 (O[19], IN1P[13], IN2);
  UB1BPPG_14_6 U15 (O[20], IN1P[14], IN2);
  UB1BPPG_15_6 U16 (O[21], IN1P[15], IN2);
  UB1BPPG_16_6 U17 (O[22], IN1P[16], IN2);
  UB1BPPG_17_6 U18 (O[23], IN1P[17], IN2);
  UB1BPPG_18_6 U19 (O[24], IN1P[18], IN2);
  UB1BPPG_19_6 U20 (O[25], IN1P[19], IN2);
  UB1BPPG_20_6 U21 (O[26], IN1P[20], IN2);
  UB1BPPG_21_6 U22 (O[27], IN1P[21], IN2);
  UB1BPPG_22_6 U23 (O[28], IN1P[22], IN2);
  UB1BPPG_23_6 U24 (O[29], IN1P[23], IN2);
  UB1BPPG_24_6 U25 (O[30], IN1P[24], IN2);
  UB1BPPG_25_6 U26 (O[31], IN1P[25], IN2);
  UB1BPPG_26_6 U27 (O[32], IN1P[26], IN2);
  UB1BPPG_27_6 U28 (O[33], IN1P[27], IN2);
  UB1BPPG_28_6 U29 (O[34], IN1P[28], IN2);
  UB1BPPG_29_6 U30 (O[35], IN1P[29], IN2);
  UB1BPPG_30_6 U31 (O[36], IN1P[30], IN2);
  NU1BPPG_31_6 U32 (NEG, IN1N, IN2);
  NUBUB1CON_37 U33 (O[37], NEG);
endmodule

module TCUVPPG_31_0_7 (O, IN1, IN2);
  output [38:7] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_7 U1 (O[7], IN1P[0], IN2);
  UB1BPPG_1_7 U2 (O[8], IN1P[1], IN2);
  UB1BPPG_2_7 U3 (O[9], IN1P[2], IN2);
  UB1BPPG_3_7 U4 (O[10], IN1P[3], IN2);
  UB1BPPG_4_7 U5 (O[11], IN1P[4], IN2);
  UB1BPPG_5_7 U6 (O[12], IN1P[5], IN2);
  UB1BPPG_6_7 U7 (O[13], IN1P[6], IN2);
  UB1BPPG_7_7 U8 (O[14], IN1P[7], IN2);
  UB1BPPG_8_7 U9 (O[15], IN1P[8], IN2);
  UB1BPPG_9_7 U10 (O[16], IN1P[9], IN2);
  UB1BPPG_10_7 U11 (O[17], IN1P[10], IN2);
  UB1BPPG_11_7 U12 (O[18], IN1P[11], IN2);
  UB1BPPG_12_7 U13 (O[19], IN1P[12], IN2);
  UB1BPPG_13_7 U14 (O[20], IN1P[13], IN2);
  UB1BPPG_14_7 U15 (O[21], IN1P[14], IN2);
  UB1BPPG_15_7 U16 (O[22], IN1P[15], IN2);
  UB1BPPG_16_7 U17 (O[23], IN1P[16], IN2);
  UB1BPPG_17_7 U18 (O[24], IN1P[17], IN2);
  UB1BPPG_18_7 U19 (O[25], IN1P[18], IN2);
  UB1BPPG_19_7 U20 (O[26], IN1P[19], IN2);
  UB1BPPG_20_7 U21 (O[27], IN1P[20], IN2);
  UB1BPPG_21_7 U22 (O[28], IN1P[21], IN2);
  UB1BPPG_22_7 U23 (O[29], IN1P[22], IN2);
  UB1BPPG_23_7 U24 (O[30], IN1P[23], IN2);
  UB1BPPG_24_7 U25 (O[31], IN1P[24], IN2);
  UB1BPPG_25_7 U26 (O[32], IN1P[25], IN2);
  UB1BPPG_26_7 U27 (O[33], IN1P[26], IN2);
  UB1BPPG_27_7 U28 (O[34], IN1P[27], IN2);
  UB1BPPG_28_7 U29 (O[35], IN1P[28], IN2);
  UB1BPPG_29_7 U30 (O[36], IN1P[29], IN2);
  UB1BPPG_30_7 U31 (O[37], IN1P[30], IN2);
  NU1BPPG_31_7 U32 (NEG, IN1N, IN2);
  NUBUB1CON_38 U33 (O[38], NEG);
endmodule

module TCUVPPG_31_0_8 (O, IN1, IN2);
  output [39:8] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_8 U1 (O[8], IN1P[0], IN2);
  UB1BPPG_1_8 U2 (O[9], IN1P[1], IN2);
  UB1BPPG_2_8 U3 (O[10], IN1P[2], IN2);
  UB1BPPG_3_8 U4 (O[11], IN1P[3], IN2);
  UB1BPPG_4_8 U5 (O[12], IN1P[4], IN2);
  UB1BPPG_5_8 U6 (O[13], IN1P[5], IN2);
  UB1BPPG_6_8 U7 (O[14], IN1P[6], IN2);
  UB1BPPG_7_8 U8 (O[15], IN1P[7], IN2);
  UB1BPPG_8_8 U9 (O[16], IN1P[8], IN2);
  UB1BPPG_9_8 U10 (O[17], IN1P[9], IN2);
  UB1BPPG_10_8 U11 (O[18], IN1P[10], IN2);
  UB1BPPG_11_8 U12 (O[19], IN1P[11], IN2);
  UB1BPPG_12_8 U13 (O[20], IN1P[12], IN2);
  UB1BPPG_13_8 U14 (O[21], IN1P[13], IN2);
  UB1BPPG_14_8 U15 (O[22], IN1P[14], IN2);
  UB1BPPG_15_8 U16 (O[23], IN1P[15], IN2);
  UB1BPPG_16_8 U17 (O[24], IN1P[16], IN2);
  UB1BPPG_17_8 U18 (O[25], IN1P[17], IN2);
  UB1BPPG_18_8 U19 (O[26], IN1P[18], IN2);
  UB1BPPG_19_8 U20 (O[27], IN1P[19], IN2);
  UB1BPPG_20_8 U21 (O[28], IN1P[20], IN2);
  UB1BPPG_21_8 U22 (O[29], IN1P[21], IN2);
  UB1BPPG_22_8 U23 (O[30], IN1P[22], IN2);
  UB1BPPG_23_8 U24 (O[31], IN1P[23], IN2);
  UB1BPPG_24_8 U25 (O[32], IN1P[24], IN2);
  UB1BPPG_25_8 U26 (O[33], IN1P[25], IN2);
  UB1BPPG_26_8 U27 (O[34], IN1P[26], IN2);
  UB1BPPG_27_8 U28 (O[35], IN1P[27], IN2);
  UB1BPPG_28_8 U29 (O[36], IN1P[28], IN2);
  UB1BPPG_29_8 U30 (O[37], IN1P[29], IN2);
  UB1BPPG_30_8 U31 (O[38], IN1P[30], IN2);
  NU1BPPG_31_8 U32 (NEG, IN1N, IN2);
  NUBUB1CON_39 U33 (O[39], NEG);
endmodule

module TCUVPPG_31_0_9 (O, IN1, IN2);
  output [40:9] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_9 U1 (O[9], IN1P[0], IN2);
  UB1BPPG_1_9 U2 (O[10], IN1P[1], IN2);
  UB1BPPG_2_9 U3 (O[11], IN1P[2], IN2);
  UB1BPPG_3_9 U4 (O[12], IN1P[3], IN2);
  UB1BPPG_4_9 U5 (O[13], IN1P[4], IN2);
  UB1BPPG_5_9 U6 (O[14], IN1P[5], IN2);
  UB1BPPG_6_9 U7 (O[15], IN1P[6], IN2);
  UB1BPPG_7_9 U8 (O[16], IN1P[7], IN2);
  UB1BPPG_8_9 U9 (O[17], IN1P[8], IN2);
  UB1BPPG_9_9 U10 (O[18], IN1P[9], IN2);
  UB1BPPG_10_9 U11 (O[19], IN1P[10], IN2);
  UB1BPPG_11_9 U12 (O[20], IN1P[11], IN2);
  UB1BPPG_12_9 U13 (O[21], IN1P[12], IN2);
  UB1BPPG_13_9 U14 (O[22], IN1P[13], IN2);
  UB1BPPG_14_9 U15 (O[23], IN1P[14], IN2);
  UB1BPPG_15_9 U16 (O[24], IN1P[15], IN2);
  UB1BPPG_16_9 U17 (O[25], IN1P[16], IN2);
  UB1BPPG_17_9 U18 (O[26], IN1P[17], IN2);
  UB1BPPG_18_9 U19 (O[27], IN1P[18], IN2);
  UB1BPPG_19_9 U20 (O[28], IN1P[19], IN2);
  UB1BPPG_20_9 U21 (O[29], IN1P[20], IN2);
  UB1BPPG_21_9 U22 (O[30], IN1P[21], IN2);
  UB1BPPG_22_9 U23 (O[31], IN1P[22], IN2);
  UB1BPPG_23_9 U24 (O[32], IN1P[23], IN2);
  UB1BPPG_24_9 U25 (O[33], IN1P[24], IN2);
  UB1BPPG_25_9 U26 (O[34], IN1P[25], IN2);
  UB1BPPG_26_9 U27 (O[35], IN1P[26], IN2);
  UB1BPPG_27_9 U28 (O[36], IN1P[27], IN2);
  UB1BPPG_28_9 U29 (O[37], IN1P[28], IN2);
  UB1BPPG_29_9 U30 (O[38], IN1P[29], IN2);
  UB1BPPG_30_9 U31 (O[39], IN1P[30], IN2);
  NU1BPPG_31_9 U32 (NEG, IN1N, IN2);
  NUBUB1CON_40 U33 (O[40], NEG);
endmodule

module UBCMBIN_32_32_31_000 (O, IN0, IN1);
  output [32:0] O;
  input IN0;
  input [31:0] IN1;
  UB1DCON_32 U0 (O[32], IN0);
  UBCON_31_0 U1 (O[31:0], IN1);
endmodule

module UBCON_10_9 (O, I);
  output [10:9] O;
  input [10:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
endmodule

module UBCON_12_10 (O, I);
  output [12:10] O;
  input [12:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
endmodule

module UBCON_14_13 (O, I);
  output [14:13] O;
  input [14:13] I;
  UB1DCON_13 U0 (O[13], I[13]);
  UB1DCON_14 U1 (O[14], I[14]);
endmodule

module UBCON_17_14 (O, I);
  output [17:14] O;
  input [17:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
endmodule

module UBCON_19_18 (O, I);
  output [19:18] O;
  input [19:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_23_22 (O, I);
  output [23:22] O;
  input [23:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
endmodule

module UBCON_24_19 (O, I);
  output [24:19] O;
  input [24:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
  UB1DCON_23 U4 (O[23], I[23]);
  UB1DCON_24 U5 (O[24], I[24]);
endmodule

module UBCON_26_25 (O, I);
  output [26:25] O;
  input [26:25] I;
  UB1DCON_25 U0 (O[25], I[25]);
  UB1DCON_26 U1 (O[26], I[26]);
endmodule

module UBCON_27_25 (O, I);
  output [27:25] O;
  input [27:25] I;
  UB1DCON_25 U0 (O[25], I[25]);
  UB1DCON_26 U1 (O[26], I[26]);
  UB1DCON_27 U2 (O[27], I[27]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_31_0 (O, I);
  output [31:0] O;
  input [31:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
  UB1DCON_28 U28 (O[28], I[28]);
  UB1DCON_29 U29 (O[29], I[29]);
  UB1DCON_30 U30 (O[30], I[30]);
  UB1DCON_31 U31 (O[31], I[31]);
endmodule

module UBCON_36_34 (O, I);
  output [36:34] O;
  input [36:34] I;
  UB1DCON_34 U0 (O[34], I[34]);
  UB1DCON_35 U1 (O[35], I[35]);
  UB1DCON_36 U2 (O[36], I[36]);
endmodule

module UBCON_39_37 (O, I);
  output [39:37] O;
  input [39:37] I;
  UB1DCON_37 U0 (O[37], I[37]);
  UB1DCON_38 U1 (O[38], I[38]);
  UB1DCON_39 U2 (O[39], I[39]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_43_40 (O, I);
  output [43:40] O;
  input [43:40] I;
  UB1DCON_40 U0 (O[40], I[40]);
  UB1DCON_41 U1 (O[41], I[41]);
  UB1DCON_42 U2 (O[42], I[42]);
  UB1DCON_43 U3 (O[43], I[43]);
endmodule

module UBCON_49_44 (O, I);
  output [49:44] O;
  input [49:44] I;
  UB1DCON_44 U0 (O[44], I[44]);
  UB1DCON_45 U1 (O[45], I[45]);
  UB1DCON_46 U2 (O[46], I[46]);
  UB1DCON_47 U3 (O[47], I[47]);
  UB1DCON_48 U4 (O[48], I[48]);
  UB1DCON_49 U5 (O[49], I[49]);
endmodule

module UBCON_49_47 (O, I);
  output [49:47] O;
  input [49:47] I;
  UB1DCON_47 U0 (O[47], I[47]);
  UB1DCON_48 U1 (O[48], I[48]);
  UB1DCON_49 U2 (O[49], I[49]);
endmodule

module UBCON_49_48 (O, I);
  output [49:48] O;
  input [49:48] I;
  UB1DCON_48 U0 (O[48], I[48]);
  UB1DCON_49 U1 (O[49], I[49]);
endmodule

module UBCON_4_0 (O, I);
  output [4:0] O;
  input [4:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
endmodule

module UBCON_58_50 (O, I);
  output [58:50] O;
  input [58:50] I;
  UB1DCON_50 U0 (O[50], I[50]);
  UB1DCON_51 U1 (O[51], I[51]);
  UB1DCON_52 U2 (O[52], I[52]);
  UB1DCON_53 U3 (O[53], I[53]);
  UB1DCON_54 U4 (O[54], I[54]);
  UB1DCON_55 U5 (O[55], I[55]);
  UB1DCON_56 U6 (O[56], I[56]);
  UB1DCON_57 U7 (O[57], I[57]);
  UB1DCON_58 U8 (O[58], I[58]);
endmodule

module UBCON_58_54 (O, I);
  output [58:54] O;
  input [58:54] I;
  UB1DCON_54 U0 (O[54], I[54]);
  UB1DCON_55 U1 (O[55], I[55]);
  UB1DCON_56 U2 (O[56], I[56]);
  UB1DCON_57 U3 (O[57], I[57]);
  UB1DCON_58 U4 (O[58], I[58]);
endmodule

module UBCON_58_55 (O, I);
  output [58:55] O;
  input [58:55] I;
  UB1DCON_55 U0 (O[55], I[55]);
  UB1DCON_56 U1 (O[56], I[56]);
  UB1DCON_57 U2 (O[57], I[57]);
  UB1DCON_58 U3 (O[58], I[58]);
endmodule

module UBCON_58_56 (O, I);
  output [58:56] O;
  input [58:56] I;
  UB1DCON_56 U0 (O[56], I[56]);
  UB1DCON_57 U1 (O[57], I[57]);
  UB1DCON_58 U2 (O[58], I[58]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_63_59 (O, I);
  output [63:59] O;
  input [63:59] I;
  UB1DCON_59 U0 (O[59], I[59]);
  UB1DCON_60 U1 (O[60], I[60]);
  UB1DCON_61 U2 (O[61], I[61]);
  UB1DCON_62 U3 (O[62], I[62]);
  UB1DCON_63 U4 (O[63], I[63]);
endmodule

module UBCON_63_9 (O, I);
  output [63:9] O;
  input [63:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
  UB1DCON_11 U2 (O[11], I[11]);
  UB1DCON_12 U3 (O[12], I[12]);
  UB1DCON_13 U4 (O[13], I[13]);
  UB1DCON_14 U5 (O[14], I[14]);
  UB1DCON_15 U6 (O[15], I[15]);
  UB1DCON_16 U7 (O[16], I[16]);
  UB1DCON_17 U8 (O[17], I[17]);
  UB1DCON_18 U9 (O[18], I[18]);
  UB1DCON_19 U10 (O[19], I[19]);
  UB1DCON_20 U11 (O[20], I[20]);
  UB1DCON_21 U12 (O[21], I[21]);
  UB1DCON_22 U13 (O[22], I[22]);
  UB1DCON_23 U14 (O[23], I[23]);
  UB1DCON_24 U15 (O[24], I[24]);
  UB1DCON_25 U16 (O[25], I[25]);
  UB1DCON_26 U17 (O[26], I[26]);
  UB1DCON_27 U18 (O[27], I[27]);
  UB1DCON_28 U19 (O[28], I[28]);
  UB1DCON_29 U20 (O[29], I[29]);
  UB1DCON_30 U21 (O[30], I[30]);
  UB1DCON_31 U22 (O[31], I[31]);
  UB1DCON_32 U23 (O[32], I[32]);
  UB1DCON_33 U24 (O[33], I[33]);
  UB1DCON_34 U25 (O[34], I[34]);
  UB1DCON_35 U26 (O[35], I[35]);
  UB1DCON_36 U27 (O[36], I[36]);
  UB1DCON_37 U28 (O[37], I[37]);
  UB1DCON_38 U29 (O[38], I[38]);
  UB1DCON_39 U30 (O[39], I[39]);
  UB1DCON_40 U31 (O[40], I[40]);
  UB1DCON_41 U32 (O[41], I[41]);
  UB1DCON_42 U33 (O[42], I[42]);
  UB1DCON_43 U34 (O[43], I[43]);
  UB1DCON_44 U35 (O[44], I[44]);
  UB1DCON_45 U36 (O[45], I[45]);
  UB1DCON_46 U37 (O[46], I[46]);
  UB1DCON_47 U38 (O[47], I[47]);
  UB1DCON_48 U39 (O[48], I[48]);
  UB1DCON_49 U40 (O[49], I[49]);
  UB1DCON_50 U41 (O[50], I[50]);
  UB1DCON_51 U42 (O[51], I[51]);
  UB1DCON_52 U43 (O[52], I[52]);
  UB1DCON_53 U44 (O[53], I[53]);
  UB1DCON_54 U45 (O[54], I[54]);
  UB1DCON_55 U46 (O[55], I[55]);
  UB1DCON_56 U47 (O[56], I[56]);
  UB1DCON_57 U48 (O[57], I[57]);
  UB1DCON_58 U49 (O[58], I[58]);
  UB1DCON_59 U50 (O[59], I[59]);
  UB1DCON_60 U51 (O[60], I[60]);
  UB1DCON_61 U52 (O[61], I[61]);
  UB1DCON_62 U53 (O[62], I[62]);
  UB1DCON_63 U54 (O[63], I[63]);
endmodule

module UBCON_6_0 (O, I);
  output [6:0] O;
  input [6:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
endmodule

module UBCON_7_0 (O, I);
  output [7:0] O;
  input [7:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
endmodule

module UBCON_8_0 (O, I);
  output [8:0] O;
  input [8:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
endmodule

module UBCON_8_7 (O, I);
  output [8:7] O;
  input [8:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
endmodule

module UBExtender_63_9_6000 (O, I);
  output [64:9] O;
  input [63:9] I;
  UBCON_63_9 U0 (O[63:9], I[63:9]);
  UBZero_64_64 U1 (O[64]);
endmodule

module UBKSA_64_9_63_0 (S, X, Y);
  output [65:0] S;
  input [64:9] X;
  input [63:0] Y;
  wire [64:9] Z;
  UBExtender_63_9_6000 U0 (Z[64:9], Y[63:9]);
  UBPureKSA_64_9 U1 (S[65:9], X[64:9], Z[64:9]);
  UBCON_8_0 U2 (S[8:0], Y[8:0]);
endmodule

module UBPureKSA_64_9 (S, X, Y);
  output [65:9] S;
  input [64:9] X;
  input [64:9] Y;
  wire C;
  UBPriKSA_64_9 U0 (S, X, Y, C);
  UBZero_9_9 U1 (C);
endmodule

module UBTCCONV63_65_0 (O, I);
  output [66:0] O;
  input [65:0] I;
  UBTC1CON66_0 U0 (O[0], I[0]);
  UBTC1CON66_1 U1 (O[1], I[1]);
  UBTC1CON66_2 U2 (O[2], I[2]);
  UBTC1CON66_3 U3 (O[3], I[3]);
  UBTC1CON66_4 U4 (O[4], I[4]);
  UBTC1CON66_5 U5 (O[5], I[5]);
  UBTC1CON66_6 U6 (O[6], I[6]);
  UBTC1CON66_7 U7 (O[7], I[7]);
  UBTC1CON66_8 U8 (O[8], I[8]);
  UBTC1CON66_9 U9 (O[9], I[9]);
  UBTC1CON66_10 U10 (O[10], I[10]);
  UBTC1CON66_11 U11 (O[11], I[11]);
  UBTC1CON66_12 U12 (O[12], I[12]);
  UBTC1CON66_13 U13 (O[13], I[13]);
  UBTC1CON66_14 U14 (O[14], I[14]);
  UBTC1CON66_15 U15 (O[15], I[15]);
  UBTC1CON66_16 U16 (O[16], I[16]);
  UBTC1CON66_17 U17 (O[17], I[17]);
  UBTC1CON66_18 U18 (O[18], I[18]);
  UBTC1CON66_19 U19 (O[19], I[19]);
  UBTC1CON66_20 U20 (O[20], I[20]);
  UBTC1CON66_21 U21 (O[21], I[21]);
  UBTC1CON66_22 U22 (O[22], I[22]);
  UBTC1CON66_23 U23 (O[23], I[23]);
  UBTC1CON66_24 U24 (O[24], I[24]);
  UBTC1CON66_25 U25 (O[25], I[25]);
  UBTC1CON66_26 U26 (O[26], I[26]);
  UBTC1CON66_27 U27 (O[27], I[27]);
  UBTC1CON66_28 U28 (O[28], I[28]);
  UBTC1CON66_29 U29 (O[29], I[29]);
  UBTC1CON66_30 U30 (O[30], I[30]);
  UBTC1CON66_31 U31 (O[31], I[31]);
  UBTC1CON66_32 U32 (O[32], I[32]);
  UBTC1CON66_33 U33 (O[33], I[33]);
  UBTC1CON66_34 U34 (O[34], I[34]);
  UBTC1CON66_35 U35 (O[35], I[35]);
  UBTC1CON66_36 U36 (O[36], I[36]);
  UBTC1CON66_37 U37 (O[37], I[37]);
  UBTC1CON66_38 U38 (O[38], I[38]);
  UBTC1CON66_39 U39 (O[39], I[39]);
  UBTC1CON66_40 U40 (O[40], I[40]);
  UBTC1CON66_41 U41 (O[41], I[41]);
  UBTC1CON66_42 U42 (O[42], I[42]);
  UBTC1CON66_43 U43 (O[43], I[43]);
  UBTC1CON66_44 U44 (O[44], I[44]);
  UBTC1CON66_45 U45 (O[45], I[45]);
  UBTC1CON66_46 U46 (O[46], I[46]);
  UBTC1CON66_47 U47 (O[47], I[47]);
  UBTC1CON66_48 U48 (O[48], I[48]);
  UBTC1CON66_49 U49 (O[49], I[49]);
  UBTC1CON66_50 U50 (O[50], I[50]);
  UBTC1CON66_51 U51 (O[51], I[51]);
  UBTC1CON66_52 U52 (O[52], I[52]);
  UBTC1CON66_53 U53 (O[53], I[53]);
  UBTC1CON66_54 U54 (O[54], I[54]);
  UBTC1CON66_55 U55 (O[55], I[55]);
  UBTC1CON66_56 U56 (O[56], I[56]);
  UBTC1CON66_57 U57 (O[57], I[57]);
  UBTC1CON66_58 U58 (O[58], I[58]);
  UBTC1CON66_59 U59 (O[59], I[59]);
  UBTC1CON66_60 U60 (O[60], I[60]);
  UBTC1CON66_61 U61 (O[61], I[61]);
  UBTC1CON66_62 U62 (O[62], I[62]);
  UBTCTCONV_65_63 U63 (O[66:63], I[65:63]);
endmodule

module WLCTR_32_0_32_1_3000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31);
  output [64:9] S1;
  output [63:0] S2;
  input [32:0] PP0;
  input [32:1] PP1;
  input [41:10] PP10;
  input [42:11] PP11;
  input [43:12] PP12;
  input [44:13] PP13;
  input [45:14] PP14;
  input [46:15] PP15;
  input [47:16] PP16;
  input [48:17] PP17;
  input [49:18] PP18;
  input [50:19] PP19;
  input [33:2] PP2;
  input [51:20] PP20;
  input [52:21] PP21;
  input [53:22] PP22;
  input [54:23] PP23;
  input [55:24] PP24;
  input [56:25] PP25;
  input [57:26] PP26;
  input [58:27] PP27;
  input [59:28] PP28;
  input [60:29] PP29;
  input [34:3] PP3;
  input [61:30] PP30;
  input [62:31] PP31;
  input [35:4] PP4;
  input [36:5] PP5;
  input [37:6] PP6;
  input [38:7] PP7;
  input [39:8] PP8;
  input [40:9] PP9;
  wire [33:2] IC0;
  wire [36:5] IC1;
  wire [55:24] IC10;
  wire [58:27] IC11;
  wire [61:30] IC12;
  wire [37:4] IC13;
  wire [44:10] IC14;
  wire [47:16] IC15;
  wire [53:20] IC16;
  wire [56:25] IC17;
  wire [62:29] IC18;
  wire [40:5] IC19;
  wire [39:8] IC2;
  wire [48:14] IC20;
  wire [54:21] IC21;
  wire [62:28] IC22;
  wire [44:6] IC23;
  wire [55:19] IC24;
  wire [63:29] IC25;
  wire [50:7] IC26;
  wire [63:26] IC27;
  wire [59:8] IC28;
  wire [42:11] IC3;
  wire [34:3] IC4;
  wire [40:7] IC5;
  wire [43:12] IC6;
  wire [46:15] IC7;
  wire [49:18] IC8;
  wire [52:21] IC9;
  wire [33:0] IS0;
  wire [36:3] IS1;
  wire [55:22] IS10;
  wire [58:25] IS11;
  wire [61:28] IS12;
  wire [39:0] IS13;
  wire [43:7] IS14;
  wire [49:13] IS15;
  wire [52:18] IS16;
  wire [58:22] IS17;
  wire [61:27] IS18;
  wire [43:0] IS19;
  wire [39:6] IS2;
  wire [49:10] IS20;
  wire [58:18] IS21;
  wire [62:25] IS22;
  wire [49:0] IS23;
  wire [58:14] IS24;
  wire [62:25] IS25;
  wire [58:0] IS26;
  wire [63:19] IS27;
  wire [63:0] IS28;
  wire [42:9] IS3;
  wire [36:0] IS4;
  wire [39:5] IS5;
  wire [43:9] IS6;
  wire [46:13] IS7;
  wire [49:16] IS8;
  wire [52:19] IS9;
  CSA_32_0_32_1_33_000 U0 (IC0, IS0, PP0, PP1, PP2);
  CSA_34_3_35_4_36_000 U1 (IC1, IS1, PP3, PP4, PP5);
  CSA_37_6_38_7_39_000 U2 (IC2, IS2, PP6, PP7, PP8);
  CSA_40_9_41_10_42000 U3 (IC3, IS3, PP9, PP10, PP11);
  CSA_33_0_33_2_36_000 U4 (IC4, IS4, IS0, IC0, IS1);
  CSA_36_5_39_6_39_000 U5 (IC5, IS5, IC1, IS2, IC2);
  CSA_42_9_42_11_43000 U6 (IC6, IS6, IS3, IC3, PP12);
  CSA_44_13_45_14_4000 U7 (IC7, IS7, PP13, PP14, PP15);
  CSA_47_16_48_17_4000 U8 (IC8, IS8, PP16, PP17, PP18);
  CSA_50_19_51_20_5000 U9 (IC9, IS9, PP19, PP20, PP21);
  CSA_53_22_54_23_5000 U10 (IC10, IS10, PP22, PP23, PP24);
  CSA_56_25_57_26_5000 U11 (IC11, IS11, PP25, PP26, PP27);
  CSA_59_28_60_29_6000 U12 (IC12, IS12, PP28, PP29, PP30);
  CSA_36_0_34_3_39_000 U13 (IC13, IS13, IS4, IC4, IS5);
  CSA_40_7_43_9_43_000 U14 (IC14, IS14, IC5, IS6, IC6);
  CSA_46_13_46_15_4000 U15 (IC15, IS15, IS7, IC7, IS8);
  CSA_49_18_52_19_5000 U16 (IC16, IS16, IC8, IS9, IC9);
  CSA_55_22_55_24_5000 U17 (IC17, IS17, IS10, IC10, IS11);
  CSA_58_27_61_28_6000 U18 (IC18, IS18, IC11, IS12, IC12);
  CSA_39_0_37_4_43_000 U19 (IC19, IS19, IS13, IC13, IS14);
  CSA_44_10_49_13_4000 U20 (IC20, IS20, IC14, IS15, IC15);
  CSA_52_18_53_20_5000 U21 (IC21, IS21, IS16, IC16, IS17);
  CSA_56_25_61_27_6000 U22 (IC22, IS22, IC17, IS18, IC18);
  CSA_43_0_40_5_49_000 U23 (IC23, IS23, IS19, IC19, IS20);
  CSA_48_14_58_18_5000 U24 (IC24, IS24, IC20, IS21, IC21);
  CSA_62_25_62_28_6000 U25 (IC25, IS25, IS22, IC22, PP31);
  CSA_49_0_44_6_58_000 U26 (IC26, IS26, IS23, IC23, IS24);
  CSA_55_19_62_25_6000 U27 (IC27, IS27, IC24, IS25, IC25);
  CSA_58_0_50_7_63_000 U28 (IC28, IS28, IS26, IC26, IS27);
  CSA_63_0_59_8_63_000 U29 (S1, S2, IS28, IC28, IC27);
endmodule


module acos_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000001100100100000000; // input=0.00048828125, output=1.57030804553
			11'd1: out = 32'b00000000000000001100100011100000; // input=0.00146484375, output=1.56933148252
			11'd2: out = 32'b00000000000000001100100011000000; // input=0.00244140625, output=1.56835491812
			11'd3: out = 32'b00000000000000001100100010100000; // input=0.00341796875, output=1.56737835139
			11'd4: out = 32'b00000000000000001100100010000000; // input=0.00439453125, output=1.5664017814
			11'd5: out = 32'b00000000000000001100100001100000; // input=0.00537109375, output=1.56542520722
			11'd6: out = 32'b00000000000000001100100001000000; // input=0.00634765625, output=1.56444862792
			11'd7: out = 32'b00000000000000001100100000100000; // input=0.00732421875, output=1.56347204256
			11'd8: out = 32'b00000000000000001100100000000000; // input=0.00830078125, output=1.56249545022
			11'd9: out = 32'b00000000000000001100011111100000; // input=0.00927734375, output=1.56151884996
			11'd10: out = 32'b00000000000000001100011111000000; // input=0.01025390625, output=1.56054224085
			11'd11: out = 32'b00000000000000001100011110100000; // input=0.01123046875, output=1.55956562196
			11'd12: out = 32'b00000000000000001100011110000000; // input=0.01220703125, output=1.55858899236
			11'd13: out = 32'b00000000000000001100011101100000; // input=0.01318359375, output=1.55761235111
			11'd14: out = 32'b00000000000000001100011101000000; // input=0.01416015625, output=1.55663569729
			11'd15: out = 32'b00000000000000001100011100100000; // input=0.01513671875, output=1.55565902996
			11'd16: out = 32'b00000000000000001100011100000000; // input=0.01611328125, output=1.55468234819
			11'd17: out = 32'b00000000000000001100011011100000; // input=0.01708984375, output=1.55370565105
			11'd18: out = 32'b00000000000000001100011011000000; // input=0.01806640625, output=1.5527289376
			11'd19: out = 32'b00000000000000001100011010100000; // input=0.01904296875, output=1.55175220692
			11'd20: out = 32'b00000000000000001100011010000000; // input=0.02001953125, output=1.55077545806
			11'd21: out = 32'b00000000000000001100011001100000; // input=0.02099609375, output=1.5497986901
			11'd22: out = 32'b00000000000000001100011001000000; // input=0.02197265625, output=1.5488219021
			11'd23: out = 32'b00000000000000001100011000100000; // input=0.02294921875, output=1.54784509314
			11'd24: out = 32'b00000000000000001100011000000000; // input=0.02392578125, output=1.54686826227
			11'd25: out = 32'b00000000000000001100010111100000; // input=0.02490234375, output=1.54589140856
			11'd26: out = 32'b00000000000000001100010111000000; // input=0.02587890625, output=1.54491453108
			11'd27: out = 32'b00000000000000001100010110100000; // input=0.02685546875, output=1.5439376289
			11'd28: out = 32'b00000000000000001100010110000000; // input=0.02783203125, output=1.54296070107
			11'd29: out = 32'b00000000000000001100010101100000; // input=0.02880859375, output=1.54198374668
			11'd30: out = 32'b00000000000000001100010101000000; // input=0.02978515625, output=1.54100676477
			11'd31: out = 32'b00000000000000001100010100100000; // input=0.03076171875, output=1.54002975443
			11'd32: out = 32'b00000000000000001100010100000000; // input=0.03173828125, output=1.5390527147
			11'd33: out = 32'b00000000000000001100010011100000; // input=0.03271484375, output=1.53807564466
			11'd34: out = 32'b00000000000000001100010011000000; // input=0.03369140625, output=1.53709854337
			11'd35: out = 32'b00000000000000001100010010100000; // input=0.03466796875, output=1.5361214099
			11'd36: out = 32'b00000000000000001100010010000000; // input=0.03564453125, output=1.5351442433
			11'd37: out = 32'b00000000000000001100010001100000; // input=0.03662109375, output=1.53416704265
			11'd38: out = 32'b00000000000000001100010001000000; // input=0.03759765625, output=1.533189807
			11'd39: out = 32'b00000000000000001100010000100000; // input=0.03857421875, output=1.53221253542
			11'd40: out = 32'b00000000000000001100010000000000; // input=0.03955078125, output=1.53123522697
			11'd41: out = 32'b00000000000000001100001111011111; // input=0.04052734375, output=1.53025788071
			11'd42: out = 32'b00000000000000001100001110111111; // input=0.04150390625, output=1.52928049571
			11'd43: out = 32'b00000000000000001100001110011111; // input=0.04248046875, output=1.52830307102
			11'd44: out = 32'b00000000000000001100001101111111; // input=0.04345703125, output=1.52732560571
			11'd45: out = 32'b00000000000000001100001101011111; // input=0.04443359375, output=1.52634809884
			11'd46: out = 32'b00000000000000001100001100111111; // input=0.04541015625, output=1.52537054947
			11'd47: out = 32'b00000000000000001100001100011111; // input=0.04638671875, output=1.52439295665
			11'd48: out = 32'b00000000000000001100001011111111; // input=0.04736328125, output=1.52341531946
			11'd49: out = 32'b00000000000000001100001011011111; // input=0.04833984375, output=1.52243763694
			11'd50: out = 32'b00000000000000001100001010111111; // input=0.04931640625, output=1.52145990816
			11'd51: out = 32'b00000000000000001100001010011111; // input=0.05029296875, output=1.52048213218
			11'd52: out = 32'b00000000000000001100001001111111; // input=0.05126953125, output=1.51950430805
			11'd53: out = 32'b00000000000000001100001001011111; // input=0.05224609375, output=1.51852643484
			11'd54: out = 32'b00000000000000001100001000111111; // input=0.05322265625, output=1.51754851159
			11'd55: out = 32'b00000000000000001100001000011111; // input=0.05419921875, output=1.51657053737
			11'd56: out = 32'b00000000000000001100000111111111; // input=0.05517578125, output=1.51559251124
			11'd57: out = 32'b00000000000000001100000111011111; // input=0.05615234375, output=1.51461443224
			11'd58: out = 32'b00000000000000001100000110111111; // input=0.05712890625, output=1.51363629943
			11'd59: out = 32'b00000000000000001100000110011111; // input=0.05810546875, output=1.51265811188
			11'd60: out = 32'b00000000000000001100000101111111; // input=0.05908203125, output=1.51167986863
			11'd61: out = 32'b00000000000000001100000101011111; // input=0.06005859375, output=1.51070156874
			11'd62: out = 32'b00000000000000001100000100111111; // input=0.06103515625, output=1.50972321126
			11'd63: out = 32'b00000000000000001100000100011111; // input=0.06201171875, output=1.50874479525
			11'd64: out = 32'b00000000000000001100000011111110; // input=0.06298828125, output=1.50776631976
			11'd65: out = 32'b00000000000000001100000011011110; // input=0.06396484375, output=1.50678778383
			11'd66: out = 32'b00000000000000001100000010111110; // input=0.06494140625, output=1.50580918653
			11'd67: out = 32'b00000000000000001100000010011110; // input=0.06591796875, output=1.5048305269
			11'd68: out = 32'b00000000000000001100000001111110; // input=0.06689453125, output=1.503851804
			11'd69: out = 32'b00000000000000001100000001011110; // input=0.06787109375, output=1.50287301687
			11'd70: out = 32'b00000000000000001100000000111110; // input=0.06884765625, output=1.50189416456
			11'd71: out = 32'b00000000000000001100000000011110; // input=0.06982421875, output=1.50091524612
			11'd72: out = 32'b00000000000000001011111111111110; // input=0.07080078125, output=1.49993626061
			11'd73: out = 32'b00000000000000001011111111011110; // input=0.07177734375, output=1.49895720706
			11'd74: out = 32'b00000000000000001011111110111110; // input=0.07275390625, output=1.49797808453
			11'd75: out = 32'b00000000000000001011111110011110; // input=0.07373046875, output=1.49699889206
			11'd76: out = 32'b00000000000000001011111101111110; // input=0.07470703125, output=1.49601962869
			11'd77: out = 32'b00000000000000001011111101011101; // input=0.07568359375, output=1.49504029348
			11'd78: out = 32'b00000000000000001011111100111101; // input=0.07666015625, output=1.49406088547
			11'd79: out = 32'b00000000000000001011111100011101; // input=0.07763671875, output=1.4930814037
			11'd80: out = 32'b00000000000000001011111011111101; // input=0.07861328125, output=1.49210184722
			11'd81: out = 32'b00000000000000001011111011011101; // input=0.07958984375, output=1.49112221506
			11'd82: out = 32'b00000000000000001011111010111101; // input=0.08056640625, output=1.49014250628
			11'd83: out = 32'b00000000000000001011111010011101; // input=0.08154296875, output=1.4891627199
			11'd84: out = 32'b00000000000000001011111001111101; // input=0.08251953125, output=1.48818285498
			11'd85: out = 32'b00000000000000001011111001011101; // input=0.08349609375, output=1.48720291055
			11'd86: out = 32'b00000000000000001011111000111101; // input=0.08447265625, output=1.48622288565
			11'd87: out = 32'b00000000000000001011111000011100; // input=0.08544921875, output=1.48524277933
			11'd88: out = 32'b00000000000000001011110111111100; // input=0.08642578125, output=1.48426259061
			11'd89: out = 32'b00000000000000001011110111011100; // input=0.08740234375, output=1.48328231853
			11'd90: out = 32'b00000000000000001011110110111100; // input=0.08837890625, output=1.48230196214
			11'd91: out = 32'b00000000000000001011110110011100; // input=0.08935546875, output=1.48132152047
			11'd92: out = 32'b00000000000000001011110101111100; // input=0.09033203125, output=1.48034099255
			11'd93: out = 32'b00000000000000001011110101011100; // input=0.09130859375, output=1.47936037742
			11'd94: out = 32'b00000000000000001011110100111100; // input=0.09228515625, output=1.47837967411
			11'd95: out = 32'b00000000000000001011110100011011; // input=0.09326171875, output=1.47739888165
			11'd96: out = 32'b00000000000000001011110011111011; // input=0.09423828125, output=1.47641799908
			11'd97: out = 32'b00000000000000001011110011011011; // input=0.09521484375, output=1.47543702542
			11'd98: out = 32'b00000000000000001011110010111011; // input=0.09619140625, output=1.47445595971
			11'd99: out = 32'b00000000000000001011110010011011; // input=0.09716796875, output=1.47347480098
			11'd100: out = 32'b00000000000000001011110001111011; // input=0.09814453125, output=1.47249354825
			11'd101: out = 32'b00000000000000001011110001011011; // input=0.09912109375, output=1.47151220056
			11'd102: out = 32'b00000000000000001011110000111010; // input=0.10009765625, output=1.47053075692
			11'd103: out = 32'b00000000000000001011110000011010; // input=0.10107421875, output=1.46954921638
			11'd104: out = 32'b00000000000000001011101111111010; // input=0.10205078125, output=1.46856757794
			11'd105: out = 32'b00000000000000001011101111011010; // input=0.10302734375, output=1.46758584064
			11'd106: out = 32'b00000000000000001011101110111010; // input=0.10400390625, output=1.4666040035
			11'd107: out = 32'b00000000000000001011101110011010; // input=0.10498046875, output=1.46562206555
			11'd108: out = 32'b00000000000000001011101101111001; // input=0.10595703125, output=1.4646400258
			11'd109: out = 32'b00000000000000001011101101011001; // input=0.10693359375, output=1.46365788327
			11'd110: out = 32'b00000000000000001011101100111001; // input=0.10791015625, output=1.46267563699
			11'd111: out = 32'b00000000000000001011101100011001; // input=0.10888671875, output=1.46169328597
			11'd112: out = 32'b00000000000000001011101011111001; // input=0.10986328125, output=1.46071082924
			11'd113: out = 32'b00000000000000001011101011011000; // input=0.11083984375, output=1.45972826581
			11'd114: out = 32'b00000000000000001011101010111000; // input=0.11181640625, output=1.45874559469
			11'd115: out = 32'b00000000000000001011101010011000; // input=0.11279296875, output=1.45776281491
			11'd116: out = 32'b00000000000000001011101001111000; // input=0.11376953125, output=1.45677992547
			11'd117: out = 32'b00000000000000001011101001011000; // input=0.11474609375, output=1.45579692539
			11'd118: out = 32'b00000000000000001011101000110111; // input=0.11572265625, output=1.45481381369
			11'd119: out = 32'b00000000000000001011101000010111; // input=0.11669921875, output=1.45383058936
			11'd120: out = 32'b00000000000000001011100111110111; // input=0.11767578125, output=1.45284725144
			11'd121: out = 32'b00000000000000001011100111010111; // input=0.11865234375, output=1.45186379891
			11'd122: out = 32'b00000000000000001011100110110110; // input=0.11962890625, output=1.4508802308
			11'd123: out = 32'b00000000000000001011100110010110; // input=0.12060546875, output=1.4498965461
			11'd124: out = 32'b00000000000000001011100101110110; // input=0.12158203125, output=1.44891274383
			11'd125: out = 32'b00000000000000001011100101010110; // input=0.12255859375, output=1.447928823
			11'd126: out = 32'b00000000000000001011100100110101; // input=0.12353515625, output=1.4469447826
			11'd127: out = 32'b00000000000000001011100100010101; // input=0.12451171875, output=1.44596062163
			11'd128: out = 32'b00000000000000001011100011110101; // input=0.12548828125, output=1.44497633911
			11'd129: out = 32'b00000000000000001011100011010101; // input=0.12646484375, output=1.44399193403
			11'd130: out = 32'b00000000000000001011100010110100; // input=0.12744140625, output=1.44300740539
			11'd131: out = 32'b00000000000000001011100010010100; // input=0.12841796875, output=1.44202275218
			11'd132: out = 32'b00000000000000001011100001110100; // input=0.12939453125, output=1.44103797342
			11'd133: out = 32'b00000000000000001011100001010100; // input=0.13037109375, output=1.44005306809
			11'd134: out = 32'b00000000000000001011100000110011; // input=0.13134765625, output=1.4390680352
			11'd135: out = 32'b00000000000000001011100000010011; // input=0.13232421875, output=1.43808287372
			11'd136: out = 32'b00000000000000001011011111110011; // input=0.13330078125, output=1.43709758266
			11'd137: out = 32'b00000000000000001011011111010011; // input=0.13427734375, output=1.43611216102
			11'd138: out = 32'b00000000000000001011011110110010; // input=0.13525390625, output=1.43512660777
			11'd139: out = 32'b00000000000000001011011110010010; // input=0.13623046875, output=1.43414092191
			11'd140: out = 32'b00000000000000001011011101110010; // input=0.13720703125, output=1.43315510243
			11'd141: out = 32'b00000000000000001011011101010001; // input=0.13818359375, output=1.43216914831
			11'd142: out = 32'b00000000000000001011011100110001; // input=0.13916015625, output=1.43118305855
			11'd143: out = 32'b00000000000000001011011100010001; // input=0.14013671875, output=1.43019683212
			11'd144: out = 32'b00000000000000001011011011110000; // input=0.14111328125, output=1.42921046801
			11'd145: out = 32'b00000000000000001011011011010000; // input=0.14208984375, output=1.4282239652
			11'd146: out = 32'b00000000000000001011011010110000; // input=0.14306640625, output=1.42723732268
			11'd147: out = 32'b00000000000000001011011010001111; // input=0.14404296875, output=1.42625053942
			11'd148: out = 32'b00000000000000001011011001101111; // input=0.14501953125, output=1.42526361439
			11'd149: out = 32'b00000000000000001011011001001111; // input=0.14599609375, output=1.42427654659
			11'd150: out = 32'b00000000000000001011011000101110; // input=0.14697265625, output=1.42328933498
			11'd151: out = 32'b00000000000000001011011000001110; // input=0.14794921875, output=1.42230197854
			11'd152: out = 32'b00000000000000001011010111101110; // input=0.14892578125, output=1.42131447624
			11'd153: out = 32'b00000000000000001011010111001101; // input=0.14990234375, output=1.42032682706
			11'd154: out = 32'b00000000000000001011010110101101; // input=0.15087890625, output=1.41933902995
			11'd155: out = 32'b00000000000000001011010110001101; // input=0.15185546875, output=1.41835108391
			11'd156: out = 32'b00000000000000001011010101101100; // input=0.15283203125, output=1.41736298788
			11'd157: out = 32'b00000000000000001011010101001100; // input=0.15380859375, output=1.41637474084
			11'd158: out = 32'b00000000000000001011010100101011; // input=0.15478515625, output=1.41538634176
			11'd159: out = 32'b00000000000000001011010100001011; // input=0.15576171875, output=1.41439778959
			11'd160: out = 32'b00000000000000001011010011101011; // input=0.15673828125, output=1.4134090833
			11'd161: out = 32'b00000000000000001011010011001010; // input=0.15771484375, output=1.41242022185
			11'd162: out = 32'b00000000000000001011010010101010; // input=0.15869140625, output=1.4114312042
			11'd163: out = 32'b00000000000000001011010010001001; // input=0.15966796875, output=1.41044202931
			11'd164: out = 32'b00000000000000001011010001101001; // input=0.16064453125, output=1.40945269613
			11'd165: out = 32'b00000000000000001011010001001001; // input=0.16162109375, output=1.40846320363
			11'd166: out = 32'b00000000000000001011010000101000; // input=0.16259765625, output=1.40747355074
			11'd167: out = 32'b00000000000000001011010000001000; // input=0.16357421875, output=1.40648373644
			11'd168: out = 32'b00000000000000001011001111100111; // input=0.16455078125, output=1.40549375965
			11'd169: out = 32'b00000000000000001011001111000111; // input=0.16552734375, output=1.40450361935
			11'd170: out = 32'b00000000000000001011001110100110; // input=0.16650390625, output=1.40351331446
			11'd171: out = 32'b00000000000000001011001110000110; // input=0.16748046875, output=1.40252284395
			11'd172: out = 32'b00000000000000001011001101100101; // input=0.16845703125, output=1.40153220675
			11'd173: out = 32'b00000000000000001011001101000101; // input=0.16943359375, output=1.40054140181
			11'd174: out = 32'b00000000000000001011001100100100; // input=0.17041015625, output=1.39955042807
			11'd175: out = 32'b00000000000000001011001100000100; // input=0.17138671875, output=1.39855928446
			11'd176: out = 32'b00000000000000001011001011100100; // input=0.17236328125, output=1.39756796994
			11'd177: out = 32'b00000000000000001011001011000011; // input=0.17333984375, output=1.39657648342
			11'd178: out = 32'b00000000000000001011001010100011; // input=0.17431640625, output=1.39558482386
			11'd179: out = 32'b00000000000000001011001010000010; // input=0.17529296875, output=1.39459299018
			11'd180: out = 32'b00000000000000001011001001100010; // input=0.17626953125, output=1.39360098132
			11'd181: out = 32'b00000000000000001011001001000001; // input=0.17724609375, output=1.3926087962
			11'd182: out = 32'b00000000000000001011001000100000; // input=0.17822265625, output=1.39161643376
			11'd183: out = 32'b00000000000000001011001000000000; // input=0.17919921875, output=1.39062389291
			11'd184: out = 32'b00000000000000001011000111011111; // input=0.18017578125, output=1.3896311726
			11'd185: out = 32'b00000000000000001011000110111111; // input=0.18115234375, output=1.38863827173
			11'd186: out = 32'b00000000000000001011000110011110; // input=0.18212890625, output=1.38764518924
			11'd187: out = 32'b00000000000000001011000101111110; // input=0.18310546875, output=1.38665192404
			11'd188: out = 32'b00000000000000001011000101011101; // input=0.18408203125, output=1.38565847506
			11'd189: out = 32'b00000000000000001011000100111101; // input=0.18505859375, output=1.3846648412
			11'd190: out = 32'b00000000000000001011000100011100; // input=0.18603515625, output=1.38367102139
			11'd191: out = 32'b00000000000000001011000011111100; // input=0.18701171875, output=1.38267701453
			11'd192: out = 32'b00000000000000001011000011011011; // input=0.18798828125, output=1.38168281954
			11'd193: out = 32'b00000000000000001011000010111010; // input=0.18896484375, output=1.38068843533
			11'd194: out = 32'b00000000000000001011000010011010; // input=0.18994140625, output=1.37969386081
			11'd195: out = 32'b00000000000000001011000001111001; // input=0.19091796875, output=1.37869909488
			11'd196: out = 32'b00000000000000001011000001011001; // input=0.19189453125, output=1.37770413645
			11'd197: out = 32'b00000000000000001011000000111000; // input=0.19287109375, output=1.37670898442
			11'd198: out = 32'b00000000000000001011000000010111; // input=0.19384765625, output=1.37571363769
			11'd199: out = 32'b00000000000000001010111111110111; // input=0.19482421875, output=1.37471809517
			11'd200: out = 32'b00000000000000001010111111010110; // input=0.19580078125, output=1.37372235573
			11'd201: out = 32'b00000000000000001010111110110101; // input=0.19677734375, output=1.3727264183
			11'd202: out = 32'b00000000000000001010111110010101; // input=0.19775390625, output=1.37173028174
			11'd203: out = 32'b00000000000000001010111101110100; // input=0.19873046875, output=1.37073394497
			11'd204: out = 32'b00000000000000001010111101010100; // input=0.19970703125, output=1.36973740686
			11'd205: out = 32'b00000000000000001010111100110011; // input=0.20068359375, output=1.36874066631
			11'd206: out = 32'b00000000000000001010111100010010; // input=0.20166015625, output=1.3677437222
			11'd207: out = 32'b00000000000000001010111011110010; // input=0.20263671875, output=1.36674657341
			11'd208: out = 32'b00000000000000001010111011010001; // input=0.20361328125, output=1.36574921883
			11'd209: out = 32'b00000000000000001010111010110000; // input=0.20458984375, output=1.36475165733
			11'd210: out = 32'b00000000000000001010111010001111; // input=0.20556640625, output=1.3637538878
			11'd211: out = 32'b00000000000000001010111001101111; // input=0.20654296875, output=1.36275590911
			11'd212: out = 32'b00000000000000001010111001001110; // input=0.20751953125, output=1.36175772013
			11'd213: out = 32'b00000000000000001010111000101101; // input=0.20849609375, output=1.36075931974
			11'd214: out = 32'b00000000000000001010111000001101; // input=0.20947265625, output=1.3597607068
			11'd215: out = 32'b00000000000000001010110111101100; // input=0.21044921875, output=1.35876188018
			11'd216: out = 32'b00000000000000001010110111001011; // input=0.21142578125, output=1.35776283875
			11'd217: out = 32'b00000000000000001010110110101010; // input=0.21240234375, output=1.35676358138
			11'd218: out = 32'b00000000000000001010110110001010; // input=0.21337890625, output=1.35576410692
			11'd219: out = 32'b00000000000000001010110101101001; // input=0.21435546875, output=1.35476441423
			11'd220: out = 32'b00000000000000001010110101001000; // input=0.21533203125, output=1.35376450217
			11'd221: out = 32'b00000000000000001010110100100111; // input=0.21630859375, output=1.35276436959
			11'd222: out = 32'b00000000000000001010110100000111; // input=0.21728515625, output=1.35176401536
			11'd223: out = 32'b00000000000000001010110011100110; // input=0.21826171875, output=1.35076343831
			11'd224: out = 32'b00000000000000001010110011000101; // input=0.21923828125, output=1.3497626373
			11'd225: out = 32'b00000000000000001010110010100100; // input=0.22021484375, output=1.34876161118
			11'd226: out = 32'b00000000000000001010110010000011; // input=0.22119140625, output=1.34776035878
			11'd227: out = 32'b00000000000000001010110001100011; // input=0.22216796875, output=1.34675887895
			11'd228: out = 32'b00000000000000001010110001000010; // input=0.22314453125, output=1.34575717054
			11'd229: out = 32'b00000000000000001010110000100001; // input=0.22412109375, output=1.34475523237
			11'd230: out = 32'b00000000000000001010110000000000; // input=0.22509765625, output=1.34375306328
			11'd231: out = 32'b00000000000000001010101111011111; // input=0.22607421875, output=1.34275066211
			11'd232: out = 32'b00000000000000001010101110111110; // input=0.22705078125, output=1.34174802769
			11'd233: out = 32'b00000000000000001010101110011110; // input=0.22802734375, output=1.34074515885
			11'd234: out = 32'b00000000000000001010101101111101; // input=0.22900390625, output=1.3397420544
			11'd235: out = 32'b00000000000000001010101101011100; // input=0.22998046875, output=1.33873871318
			11'd236: out = 32'b00000000000000001010101100111011; // input=0.23095703125, output=1.33773513401
			11'd237: out = 32'b00000000000000001010101100011010; // input=0.23193359375, output=1.3367313157
			11'd238: out = 32'b00000000000000001010101011111001; // input=0.23291015625, output=1.33572725708
			11'd239: out = 32'b00000000000000001010101011011000; // input=0.23388671875, output=1.33472295695
			11'd240: out = 32'b00000000000000001010101010110111; // input=0.23486328125, output=1.33371841413
			11'd241: out = 32'b00000000000000001010101010010110; // input=0.23583984375, output=1.33271362743
			11'd242: out = 32'b00000000000000001010101001110101; // input=0.23681640625, output=1.33170859566
			11'd243: out = 32'b00000000000000001010101001010100; // input=0.23779296875, output=1.33070331761
			11'd244: out = 32'b00000000000000001010101000110100; // input=0.23876953125, output=1.3296977921
			11'd245: out = 32'b00000000000000001010101000010011; // input=0.23974609375, output=1.32869201792
			11'd246: out = 32'b00000000000000001010100111110010; // input=0.24072265625, output=1.32768599387
			11'd247: out = 32'b00000000000000001010100111010001; // input=0.24169921875, output=1.32667971875
			11'd248: out = 32'b00000000000000001010100110110000; // input=0.24267578125, output=1.32567319134
			11'd249: out = 32'b00000000000000001010100110001111; // input=0.24365234375, output=1.32466641044
			11'd250: out = 32'b00000000000000001010100101101110; // input=0.24462890625, output=1.32365937483
			11'd251: out = 32'b00000000000000001010100101001101; // input=0.24560546875, output=1.3226520833
			11'd252: out = 32'b00000000000000001010100100101100; // input=0.24658203125, output=1.32164453463
			11'd253: out = 32'b00000000000000001010100100001011; // input=0.24755859375, output=1.3206367276
			11'd254: out = 32'b00000000000000001010100011101010; // input=0.24853515625, output=1.31962866098
			11'd255: out = 32'b00000000000000001010100011001001; // input=0.24951171875, output=1.31862033355
			11'd256: out = 32'b00000000000000001010100010101000; // input=0.25048828125, output=1.31761174409
			11'd257: out = 32'b00000000000000001010100010000110; // input=0.25146484375, output=1.31660289135
			11'd258: out = 32'b00000000000000001010100001100101; // input=0.25244140625, output=1.31559377412
			11'd259: out = 32'b00000000000000001010100001000100; // input=0.25341796875, output=1.31458439114
			11'd260: out = 32'b00000000000000001010100000100011; // input=0.25439453125, output=1.31357474118
			11'd261: out = 32'b00000000000000001010100000000010; // input=0.25537109375, output=1.312564823
			11'd262: out = 32'b00000000000000001010011111100001; // input=0.25634765625, output=1.31155463536
			11'd263: out = 32'b00000000000000001010011111000000; // input=0.25732421875, output=1.310544177
			11'd264: out = 32'b00000000000000001010011110011111; // input=0.25830078125, output=1.30953344668
			11'd265: out = 32'b00000000000000001010011101111110; // input=0.25927734375, output=1.30852244314
			11'd266: out = 32'b00000000000000001010011101011101; // input=0.26025390625, output=1.30751116513
			11'd267: out = 32'b00000000000000001010011100111011; // input=0.26123046875, output=1.30649961139
			11'd268: out = 32'b00000000000000001010011100011010; // input=0.26220703125, output=1.30548778065
			11'd269: out = 32'b00000000000000001010011011111001; // input=0.26318359375, output=1.30447567165
			11'd270: out = 32'b00000000000000001010011011011000; // input=0.26416015625, output=1.30346328313
			11'd271: out = 32'b00000000000000001010011010110111; // input=0.26513671875, output=1.30245061382
			11'd272: out = 32'b00000000000000001010011010010110; // input=0.26611328125, output=1.30143766244
			11'd273: out = 32'b00000000000000001010011001110100; // input=0.26708984375, output=1.30042442771
			11'd274: out = 32'b00000000000000001010011001010011; // input=0.26806640625, output=1.29941090836
			11'd275: out = 32'b00000000000000001010011000110010; // input=0.26904296875, output=1.2983971031
			11'd276: out = 32'b00000000000000001010011000010001; // input=0.27001953125, output=1.29738301066
			11'd277: out = 32'b00000000000000001010010111101111; // input=0.27099609375, output=1.29636862973
			11'd278: out = 32'b00000000000000001010010111001110; // input=0.27197265625, output=1.29535395904
			11'd279: out = 32'b00000000000000001010010110101101; // input=0.27294921875, output=1.29433899728
			11'd280: out = 32'b00000000000000001010010110001100; // input=0.27392578125, output=1.29332374316
			11'd281: out = 32'b00000000000000001010010101101010; // input=0.27490234375, output=1.29230819538
			11'd282: out = 32'b00000000000000001010010101001001; // input=0.27587890625, output=1.29129235264
			11'd283: out = 32'b00000000000000001010010100101000; // input=0.27685546875, output=1.29027621363
			11'd284: out = 32'b00000000000000001010010100000110; // input=0.27783203125, output=1.28925977704
			11'd285: out = 32'b00000000000000001010010011100101; // input=0.27880859375, output=1.28824304155
			11'd286: out = 32'b00000000000000001010010011000100; // input=0.27978515625, output=1.28722600586
			11'd287: out = 32'b00000000000000001010010010100010; // input=0.28076171875, output=1.28620866864
			11'd288: out = 32'b00000000000000001010010010000001; // input=0.28173828125, output=1.28519102857
			11'd289: out = 32'b00000000000000001010010001100000; // input=0.28271484375, output=1.28417308432
			11'd290: out = 32'b00000000000000001010010000111110; // input=0.28369140625, output=1.28315483458
			11'd291: out = 32'b00000000000000001010010000011101; // input=0.28466796875, output=1.28213627799
			11'd292: out = 32'b00000000000000001010001111111100; // input=0.28564453125, output=1.28111741324
			11'd293: out = 32'b00000000000000001010001111011010; // input=0.28662109375, output=1.28009823898
			11'd294: out = 32'b00000000000000001010001110111001; // input=0.28759765625, output=1.27907875386
			11'd295: out = 32'b00000000000000001010001110010111; // input=0.28857421875, output=1.27805895655
			11'd296: out = 32'b00000000000000001010001101110110; // input=0.28955078125, output=1.2770388457
			11'd297: out = 32'b00000000000000001010001101010101; // input=0.29052734375, output=1.27601841995
			11'd298: out = 32'b00000000000000001010001100110011; // input=0.29150390625, output=1.27499767795
			11'd299: out = 32'b00000000000000001010001100010010; // input=0.29248046875, output=1.27397661833
			11'd300: out = 32'b00000000000000001010001011110000; // input=0.29345703125, output=1.27295523974
			11'd301: out = 32'b00000000000000001010001011001111; // input=0.29443359375, output=1.27193354082
			11'd302: out = 32'b00000000000000001010001010101101; // input=0.29541015625, output=1.27091152019
			11'd303: out = 32'b00000000000000001010001010001100; // input=0.29638671875, output=1.26988917647
			11'd304: out = 32'b00000000000000001010001001101010; // input=0.29736328125, output=1.2688665083
			11'd305: out = 32'b00000000000000001010001001001001; // input=0.29833984375, output=1.2678435143
			11'd306: out = 32'b00000000000000001010001000100111; // input=0.29931640625, output=1.26682019307
			11'd307: out = 32'b00000000000000001010001000000110; // input=0.30029296875, output=1.26579654324
			11'd308: out = 32'b00000000000000001010000111100100; // input=0.30126953125, output=1.26477256342
			11'd309: out = 32'b00000000000000001010000111000011; // input=0.30224609375, output=1.2637482522
			11'd310: out = 32'b00000000000000001010000110100001; // input=0.30322265625, output=1.26272360819
			11'd311: out = 32'b00000000000000001010000101111111; // input=0.30419921875, output=1.26169863
			11'd312: out = 32'b00000000000000001010000101011110; // input=0.30517578125, output=1.2606733162
			11'd313: out = 32'b00000000000000001010000100111100; // input=0.30615234375, output=1.25964766541
			11'd314: out = 32'b00000000000000001010000100011011; // input=0.30712890625, output=1.2586216762
			11'd315: out = 32'b00000000000000001010000011111001; // input=0.30810546875, output=1.25759534715
			11'd316: out = 32'b00000000000000001010000011010111; // input=0.30908203125, output=1.25656867686
			11'd317: out = 32'b00000000000000001010000010110110; // input=0.31005859375, output=1.25554166389
			11'd318: out = 32'b00000000000000001010000010010100; // input=0.31103515625, output=1.25451430681
			11'd319: out = 32'b00000000000000001010000001110010; // input=0.31201171875, output=1.2534866042
			11'd320: out = 32'b00000000000000001010000001010001; // input=0.31298828125, output=1.25245855461
			11'd321: out = 32'b00000000000000001010000000101111; // input=0.31396484375, output=1.25143015662
			11'd322: out = 32'b00000000000000001010000000001101; // input=0.31494140625, output=1.25040140877
			11'd323: out = 32'b00000000000000001001111111101011; // input=0.31591796875, output=1.24937230962
			11'd324: out = 32'b00000000000000001001111111001010; // input=0.31689453125, output=1.24834285773
			11'd325: out = 32'b00000000000000001001111110101000; // input=0.31787109375, output=1.24731305162
			11'd326: out = 32'b00000000000000001001111110000110; // input=0.31884765625, output=1.24628288985
			11'd327: out = 32'b00000000000000001001111101100100; // input=0.31982421875, output=1.24525237094
			11'd328: out = 32'b00000000000000001001111101000011; // input=0.32080078125, output=1.24422149344
			11'd329: out = 32'b00000000000000001001111100100001; // input=0.32177734375, output=1.24319025588
			11'd330: out = 32'b00000000000000001001111011111111; // input=0.32275390625, output=1.24215865677
			11'd331: out = 32'b00000000000000001001111011011101; // input=0.32373046875, output=1.24112669464
			11'd332: out = 32'b00000000000000001001111010111011; // input=0.32470703125, output=1.240094368
			11'd333: out = 32'b00000000000000001001111010011010; // input=0.32568359375, output=1.23906167537
			11'd334: out = 32'b00000000000000001001111001111000; // input=0.32666015625, output=1.23802861525
			11'd335: out = 32'b00000000000000001001111001010110; // input=0.32763671875, output=1.23699518615
			11'd336: out = 32'b00000000000000001001111000110100; // input=0.32861328125, output=1.23596138656
			11'd337: out = 32'b00000000000000001001111000010010; // input=0.32958984375, output=1.23492721499
			11'd338: out = 32'b00000000000000001001110111110000; // input=0.33056640625, output=1.23389266992
			11'd339: out = 32'b00000000000000001001110111001110; // input=0.33154296875, output=1.23285774984
			11'd340: out = 32'b00000000000000001001110110101100; // input=0.33251953125, output=1.23182245324
			11'd341: out = 32'b00000000000000001001110110001010; // input=0.33349609375, output=1.23078677858
			11'd342: out = 32'b00000000000000001001110101101000; // input=0.33447265625, output=1.22975072435
			11'd343: out = 32'b00000000000000001001110101000111; // input=0.33544921875, output=1.228714289
			11'd344: out = 32'b00000000000000001001110100100101; // input=0.33642578125, output=1.22767747102
			11'd345: out = 32'b00000000000000001001110100000011; // input=0.33740234375, output=1.22664026885
			11'd346: out = 32'b00000000000000001001110011100001; // input=0.33837890625, output=1.22560268096
			11'd347: out = 32'b00000000000000001001110010111111; // input=0.33935546875, output=1.22456470579
			11'd348: out = 32'b00000000000000001001110010011101; // input=0.34033203125, output=1.22352634178
			11'd349: out = 32'b00000000000000001001110001111010; // input=0.34130859375, output=1.22248758739
			11'd350: out = 32'b00000000000000001001110001011000; // input=0.34228515625, output=1.22144844105
			11'd351: out = 32'b00000000000000001001110000110110; // input=0.34326171875, output=1.22040890119
			11'd352: out = 32'b00000000000000001001110000010100; // input=0.34423828125, output=1.21936896624
			11'd353: out = 32'b00000000000000001001101111110010; // input=0.34521484375, output=1.21832863463
			11'd354: out = 32'b00000000000000001001101111010000; // input=0.34619140625, output=1.21728790476
			11'd355: out = 32'b00000000000000001001101110101110; // input=0.34716796875, output=1.21624677506
			11'd356: out = 32'b00000000000000001001101110001100; // input=0.34814453125, output=1.21520524394
			11'd357: out = 32'b00000000000000001001101101101010; // input=0.34912109375, output=1.21416330979
			11'd358: out = 32'b00000000000000001001101101001000; // input=0.35009765625, output=1.21312097102
			11'd359: out = 32'b00000000000000001001101100100101; // input=0.35107421875, output=1.21207822602
			11'd360: out = 32'b00000000000000001001101100000011; // input=0.35205078125, output=1.21103507318
			11'd361: out = 32'b00000000000000001001101011100001; // input=0.35302734375, output=1.20999151089
			11'd362: out = 32'b00000000000000001001101010111111; // input=0.35400390625, output=1.20894753753
			11'd363: out = 32'b00000000000000001001101010011101; // input=0.35498046875, output=1.20790315147
			11'd364: out = 32'b00000000000000001001101001111010; // input=0.35595703125, output=1.20685835107
			11'd365: out = 32'b00000000000000001001101001011000; // input=0.35693359375, output=1.20581313471
			11'd366: out = 32'b00000000000000001001101000110110; // input=0.35791015625, output=1.20476750075
			11'd367: out = 32'b00000000000000001001101000010100; // input=0.35888671875, output=1.20372144753
			11'd368: out = 32'b00000000000000001001100111110001; // input=0.35986328125, output=1.20267497342
			11'd369: out = 32'b00000000000000001001100111001111; // input=0.36083984375, output=1.20162807674
			11'd370: out = 32'b00000000000000001001100110101101; // input=0.36181640625, output=1.20058075585
			11'd371: out = 32'b00000000000000001001100110001010; // input=0.36279296875, output=1.19953300907
			11'd372: out = 32'b00000000000000001001100101101000; // input=0.36376953125, output=1.19848483473
			11'd373: out = 32'b00000000000000001001100101000110; // input=0.36474609375, output=1.19743623116
			11'd374: out = 32'b00000000000000001001100100100011; // input=0.36572265625, output=1.19638719668
			11'd375: out = 32'b00000000000000001001100100000001; // input=0.36669921875, output=1.19533772959
			11'd376: out = 32'b00000000000000001001100011011110; // input=0.36767578125, output=1.19428782821
			11'd377: out = 32'b00000000000000001001100010111100; // input=0.36865234375, output=1.19323749083
			11'd378: out = 32'b00000000000000001001100010011010; // input=0.36962890625, output=1.19218671575
			11'd379: out = 32'b00000000000000001001100001110111; // input=0.37060546875, output=1.19113550126
			11'd380: out = 32'b00000000000000001001100001010101; // input=0.37158203125, output=1.19008384566
			11'd381: out = 32'b00000000000000001001100000110010; // input=0.37255859375, output=1.1890317472
			11'd382: out = 32'b00000000000000001001100000010000; // input=0.37353515625, output=1.18797920418
			11'd383: out = 32'b00000000000000001001011111101101; // input=0.37451171875, output=1.18692621486
			11'd384: out = 32'b00000000000000001001011111001011; // input=0.37548828125, output=1.18587277751
			11'd385: out = 32'b00000000000000001001011110101000; // input=0.37646484375, output=1.18481889037
			11'd386: out = 32'b00000000000000001001011110000110; // input=0.37744140625, output=1.1837645517
			11'd387: out = 32'b00000000000000001001011101100011; // input=0.37841796875, output=1.18270975975
			11'd388: out = 32'b00000000000000001001011101000000; // input=0.37939453125, output=1.18165451275
			11'd389: out = 32'b00000000000000001001011100011110; // input=0.38037109375, output=1.18059880895
			11'd390: out = 32'b00000000000000001001011011111011; // input=0.38134765625, output=1.17954264656
			11'd391: out = 32'b00000000000000001001011011011001; // input=0.38232421875, output=1.17848602382
			11'd392: out = 32'b00000000000000001001011010110110; // input=0.38330078125, output=1.17742893893
			11'd393: out = 32'b00000000000000001001011010010011; // input=0.38427734375, output=1.17637139011
			11'd394: out = 32'b00000000000000001001011001110001; // input=0.38525390625, output=1.17531337555
			11'd395: out = 32'b00000000000000001001011001001110; // input=0.38623046875, output=1.17425489347
			11'd396: out = 32'b00000000000000001001011000101011; // input=0.38720703125, output=1.17319594205
			11'd397: out = 32'b00000000000000001001011000001001; // input=0.38818359375, output=1.17213651948
			11'd398: out = 32'b00000000000000001001010111100110; // input=0.38916015625, output=1.17107662394
			11'd399: out = 32'b00000000000000001001010111000011; // input=0.39013671875, output=1.17001625359
			11'd400: out = 32'b00000000000000001001010110100000; // input=0.39111328125, output=1.16895540662
			11'd401: out = 32'b00000000000000001001010101111110; // input=0.39208984375, output=1.16789408118
			11'd402: out = 32'b00000000000000001001010101011011; // input=0.39306640625, output=1.16683227542
			11'd403: out = 32'b00000000000000001001010100111000; // input=0.39404296875, output=1.16576998749
			11'd404: out = 32'b00000000000000001001010100010101; // input=0.39501953125, output=1.16470721554
			11'd405: out = 32'b00000000000000001001010011110010; // input=0.39599609375, output=1.1636439577
			11'd406: out = 32'b00000000000000001001010011001111; // input=0.39697265625, output=1.16258021211
			11'd407: out = 32'b00000000000000001001010010101101; // input=0.39794921875, output=1.16151597687
			11'd408: out = 32'b00000000000000001001010010001010; // input=0.39892578125, output=1.16045125012
			11'd409: out = 32'b00000000000000001001010001100111; // input=0.39990234375, output=1.15938602995
			11'd410: out = 32'b00000000000000001001010001000100; // input=0.40087890625, output=1.15832031448
			11'd411: out = 32'b00000000000000001001010000100001; // input=0.40185546875, output=1.1572541018
			11'd412: out = 32'b00000000000000001001001111111110; // input=0.40283203125, output=1.15618738999
			11'd413: out = 32'b00000000000000001001001111011011; // input=0.40380859375, output=1.15512017715
			11'd414: out = 32'b00000000000000001001001110111000; // input=0.40478515625, output=1.15405246134
			11'd415: out = 32'b00000000000000001001001110010101; // input=0.40576171875, output=1.15298424064
			11'd416: out = 32'b00000000000000001001001101110010; // input=0.40673828125, output=1.15191551311
			11'd417: out = 32'b00000000000000001001001101001111; // input=0.40771484375, output=1.1508462768
			11'd418: out = 32'b00000000000000001001001100101100; // input=0.40869140625, output=1.14977652977
			11'd419: out = 32'b00000000000000001001001100001001; // input=0.40966796875, output=1.14870627005
			11'd420: out = 32'b00000000000000001001001011100110; // input=0.41064453125, output=1.14763549568
			11'd421: out = 32'b00000000000000001001001011000011; // input=0.41162109375, output=1.14656420469
			11'd422: out = 32'b00000000000000001001001010011111; // input=0.41259765625, output=1.14549239509
			11'd423: out = 32'b00000000000000001001001001111100; // input=0.41357421875, output=1.1444200649
			11'd424: out = 32'b00000000000000001001001001011001; // input=0.41455078125, output=1.14334721213
			11'd425: out = 32'b00000000000000001001001000110110; // input=0.41552734375, output=1.14227383477
			11'd426: out = 32'b00000000000000001001001000010011; // input=0.41650390625, output=1.14119993082
			11'd427: out = 32'b00000000000000001001000111110000; // input=0.41748046875, output=1.14012549826
			11'd428: out = 32'b00000000000000001001000111001100; // input=0.41845703125, output=1.13905053506
			11'd429: out = 32'b00000000000000001001000110101001; // input=0.41943359375, output=1.1379750392
			11'd430: out = 32'b00000000000000001001000110000110; // input=0.42041015625, output=1.13689900863
			11'd431: out = 32'b00000000000000001001000101100011; // input=0.42138671875, output=1.13582244131
			11'd432: out = 32'b00000000000000001001000100111111; // input=0.42236328125, output=1.13474533519
			11'd433: out = 32'b00000000000000001001000100011100; // input=0.42333984375, output=1.13366768821
			11'd434: out = 32'b00000000000000001001000011111001; // input=0.42431640625, output=1.13258949829
			11'd435: out = 32'b00000000000000001001000011010101; // input=0.42529296875, output=1.13151076336
			11'd436: out = 32'b00000000000000001001000010110010; // input=0.42626953125, output=1.13043148133
			11'd437: out = 32'b00000000000000001001000010001111; // input=0.42724609375, output=1.12935165012
			11'd438: out = 32'b00000000000000001001000001101011; // input=0.42822265625, output=1.12827126762
			11'd439: out = 32'b00000000000000001001000001001000; // input=0.42919921875, output=1.12719033172
			11'd440: out = 32'b00000000000000001001000000100100; // input=0.43017578125, output=1.12610884031
			11'd441: out = 32'b00000000000000001001000000000001; // input=0.43115234375, output=1.12502679127
			11'd442: out = 32'b00000000000000001000111111011101; // input=0.43212890625, output=1.12394418246
			11'd443: out = 32'b00000000000000001000111110111010; // input=0.43310546875, output=1.12286101173
			11'd444: out = 32'b00000000000000001000111110010110; // input=0.43408203125, output=1.12177727695
			11'd445: out = 32'b00000000000000001000111101110011; // input=0.43505859375, output=1.12069297596
			11'd446: out = 32'b00000000000000001000111101001111; // input=0.43603515625, output=1.11960810658
			11'd447: out = 32'b00000000000000001000111100101100; // input=0.43701171875, output=1.11852266665
			11'd448: out = 32'b00000000000000001000111100001000; // input=0.43798828125, output=1.11743665399
			11'd449: out = 32'b00000000000000001000111011100101; // input=0.43896484375, output=1.1163500664
			11'd450: out = 32'b00000000000000001000111011000001; // input=0.43994140625, output=1.11526290168
			11'd451: out = 32'b00000000000000001000111010011101; // input=0.44091796875, output=1.11417515763
			11'd452: out = 32'b00000000000000001000111001111010; // input=0.44189453125, output=1.11308683204
			11'd453: out = 32'b00000000000000001000111001010110; // input=0.44287109375, output=1.11199792267
			11'd454: out = 32'b00000000000000001000111000110010; // input=0.44384765625, output=1.11090842729
			11'd455: out = 32'b00000000000000001000111000001111; // input=0.44482421875, output=1.10981834366
			11'd456: out = 32'b00000000000000001000110111101011; // input=0.44580078125, output=1.10872766953
			11'd457: out = 32'b00000000000000001000110111000111; // input=0.44677734375, output=1.10763640264
			11'd458: out = 32'b00000000000000001000110110100011; // input=0.44775390625, output=1.10654454072
			11'd459: out = 32'b00000000000000001000110101111111; // input=0.44873046875, output=1.10545208149
			11'd460: out = 32'b00000000000000001000110101011100; // input=0.44970703125, output=1.10435902266
			11'd461: out = 32'b00000000000000001000110100111000; // input=0.45068359375, output=1.10326536194
			11'd462: out = 32'b00000000000000001000110100010100; // input=0.45166015625, output=1.10217109702
			11'd463: out = 32'b00000000000000001000110011110000; // input=0.45263671875, output=1.10107622559
			11'd464: out = 32'b00000000000000001000110011001100; // input=0.45361328125, output=1.09998074532
			11'd465: out = 32'b00000000000000001000110010101000; // input=0.45458984375, output=1.09888465389
			11'd466: out = 32'b00000000000000001000110010000100; // input=0.45556640625, output=1.09778794893
			11'd467: out = 32'b00000000000000001000110001100000; // input=0.45654296875, output=1.09669062811
			11'd468: out = 32'b00000000000000001000110000111100; // input=0.45751953125, output=1.09559268906
			11'd469: out = 32'b00000000000000001000110000011000; // input=0.45849609375, output=1.09449412941
			11'd470: out = 32'b00000000000000001000101111110100; // input=0.45947265625, output=1.09339494678
			11'd471: out = 32'b00000000000000001000101111010000; // input=0.46044921875, output=1.09229513877
			11'd472: out = 32'b00000000000000001000101110101100; // input=0.46142578125, output=1.09119470298
			11'd473: out = 32'b00000000000000001000101110001000; // input=0.46240234375, output=1.09009363702
			11'd474: out = 32'b00000000000000001000101101100100; // input=0.46337890625, output=1.08899193844
			11'd475: out = 32'b00000000000000001000101101000000; // input=0.46435546875, output=1.08788960482
			11'd476: out = 32'b00000000000000001000101100011100; // input=0.46533203125, output=1.08678663373
			11'd477: out = 32'b00000000000000001000101011111000; // input=0.46630859375, output=1.0856830227
			11'd478: out = 32'b00000000000000001000101011010011; // input=0.46728515625, output=1.08457876928
			11'd479: out = 32'b00000000000000001000101010101111; // input=0.46826171875, output=1.083473871
			11'd480: out = 32'b00000000000000001000101010001011; // input=0.46923828125, output=1.08236832536
			11'd481: out = 32'b00000000000000001000101001100111; // input=0.47021484375, output=1.08126212989
			11'd482: out = 32'b00000000000000001000101001000011; // input=0.47119140625, output=1.08015528208
			11'd483: out = 32'b00000000000000001000101000011110; // input=0.47216796875, output=1.07904777941
			11'd484: out = 32'b00000000000000001000100111111010; // input=0.47314453125, output=1.07793961935
			11'd485: out = 32'b00000000000000001000100111010110; // input=0.47412109375, output=1.07683079938
			11'd486: out = 32'b00000000000000001000100110110001; // input=0.47509765625, output=1.07572131695
			11'd487: out = 32'b00000000000000001000100110001101; // input=0.47607421875, output=1.0746111695
			11'd488: out = 32'b00000000000000001000100101101000; // input=0.47705078125, output=1.07350035446
			11'd489: out = 32'b00000000000000001000100101000100; // input=0.47802734375, output=1.07238886925
			11'd490: out = 32'b00000000000000001000100100100000; // input=0.47900390625, output=1.07127671129
			11'd491: out = 32'b00000000000000001000100011111011; // input=0.47998046875, output=1.07016387796
			11'd492: out = 32'b00000000000000001000100011010111; // input=0.48095703125, output=1.06905036667
			11'd493: out = 32'b00000000000000001000100010110010; // input=0.48193359375, output=1.06793617478
			11'd494: out = 32'b00000000000000001000100010001110; // input=0.48291015625, output=1.06682129967
			11'd495: out = 32'b00000000000000001000100001101001; // input=0.48388671875, output=1.06570573867
			11'd496: out = 32'b00000000000000001000100001000100; // input=0.48486328125, output=1.06458948915
			11'd497: out = 32'b00000000000000001000100000100000; // input=0.48583984375, output=1.06347254841
			11'd498: out = 32'b00000000000000001000011111111011; // input=0.48681640625, output=1.0623549138
			11'd499: out = 32'b00000000000000001000011111010111; // input=0.48779296875, output=1.0612365826
			11'd500: out = 32'b00000000000000001000011110110010; // input=0.48876953125, output=1.06011755212
			11'd501: out = 32'b00000000000000001000011110001101; // input=0.48974609375, output=1.05899781963
			11'd502: out = 32'b00000000000000001000011101101001; // input=0.49072265625, output=1.05787738241
			11'd503: out = 32'b00000000000000001000011101000100; // input=0.49169921875, output=1.05675623772
			11'd504: out = 32'b00000000000000001000011100011111; // input=0.49267578125, output=1.05563438281
			11'd505: out = 32'b00000000000000001000011011111010; // input=0.49365234375, output=1.0545118149
			11'd506: out = 32'b00000000000000001000011011010101; // input=0.49462890625, output=1.05338853122
			11'd507: out = 32'b00000000000000001000011010110001; // input=0.49560546875, output=1.05226452897
			11'd508: out = 32'b00000000000000001000011010001100; // input=0.49658203125, output=1.05113980536
			11'd509: out = 32'b00000000000000001000011001100111; // input=0.49755859375, output=1.05001435757
			11'd510: out = 32'b00000000000000001000011001000010; // input=0.49853515625, output=1.04888818277
			11'd511: out = 32'b00000000000000001000011000011101; // input=0.49951171875, output=1.04776127811
			11'd512: out = 32'b00000000000000001000010111111000; // input=0.50048828125, output=1.04663364075
			11'd513: out = 32'b00000000000000001000010111010011; // input=0.50146484375, output=1.04550526781
			11'd514: out = 32'b00000000000000001000010110101110; // input=0.50244140625, output=1.04437615641
			11'd515: out = 32'b00000000000000001000010110001001; // input=0.50341796875, output=1.04324630367
			11'd516: out = 32'b00000000000000001000010101100100; // input=0.50439453125, output=1.04211570666
			11'd517: out = 32'b00000000000000001000010100111111; // input=0.50537109375, output=1.04098436248
			11'd518: out = 32'b00000000000000001000010100011010; // input=0.50634765625, output=1.03985226819
			11'd519: out = 32'b00000000000000001000010011110101; // input=0.50732421875, output=1.03871942083
			11'd520: out = 32'b00000000000000001000010011010000; // input=0.50830078125, output=1.03758581745
			11'd521: out = 32'b00000000000000001000010010101010; // input=0.50927734375, output=1.03645145508
			11'd522: out = 32'b00000000000000001000010010000101; // input=0.51025390625, output=1.03531633071
			11'd523: out = 32'b00000000000000001000010001100000; // input=0.51123046875, output=1.03418044136
			11'd524: out = 32'b00000000000000001000010000111011; // input=0.51220703125, output=1.033043784
			11'd525: out = 32'b00000000000000001000010000010110; // input=0.51318359375, output=1.03190635561
			11'd526: out = 32'b00000000000000001000001111110000; // input=0.51416015625, output=1.03076815313
			11'd527: out = 32'b00000000000000001000001111001011; // input=0.51513671875, output=1.0296291735
			11'd528: out = 32'b00000000000000001000001110100110; // input=0.51611328125, output=1.02848941365
			11'd529: out = 32'b00000000000000001000001110000000; // input=0.51708984375, output=1.0273488705
			11'd530: out = 32'b00000000000000001000001101011011; // input=0.51806640625, output=1.02620754093
			11'd531: out = 32'b00000000000000001000001100110101; // input=0.51904296875, output=1.02506542184
			11'd532: out = 32'b00000000000000001000001100010000; // input=0.52001953125, output=1.02392251008
			11'd533: out = 32'b00000000000000001000001011101010; // input=0.52099609375, output=1.0227788025
			11'd534: out = 32'b00000000000000001000001011000101; // input=0.52197265625, output=1.02163429595
			11'd535: out = 32'b00000000000000001000001010011111; // input=0.52294921875, output=1.02048898724
			11'd536: out = 32'b00000000000000001000001001111010; // input=0.52392578125, output=1.01934287318
			11'd537: out = 32'b00000000000000001000001001010100; // input=0.52490234375, output=1.01819595056
			11'd538: out = 32'b00000000000000001000001000101111; // input=0.52587890625, output=1.01704821615
			11'd539: out = 32'b00000000000000001000001000001001; // input=0.52685546875, output=1.01589966671
			11'd540: out = 32'b00000000000000001000000111100011; // input=0.52783203125, output=1.01475029899
			11'd541: out = 32'b00000000000000001000000110111110; // input=0.52880859375, output=1.01360010971
			11'd542: out = 32'b00000000000000001000000110011000; // input=0.52978515625, output=1.01244909558
			11'd543: out = 32'b00000000000000001000000101110010; // input=0.53076171875, output=1.0112972533
			11'd544: out = 32'b00000000000000001000000101001100; // input=0.53173828125, output=1.01014457955
			11'd545: out = 32'b00000000000000001000000100100111; // input=0.53271484375, output=1.00899107098
			11'd546: out = 32'b00000000000000001000000100000001; // input=0.53369140625, output=1.00783672425
			11'd547: out = 32'b00000000000000001000000011011011; // input=0.53466796875, output=1.00668153598
			11'd548: out = 32'b00000000000000001000000010110101; // input=0.53564453125, output=1.00552550278
			11'd549: out = 32'b00000000000000001000000010001111; // input=0.53662109375, output=1.00436862125
			11'd550: out = 32'b00000000000000001000000001101001; // input=0.53759765625, output=1.00321088797
			11'd551: out = 32'b00000000000000001000000001000011; // input=0.53857421875, output=1.00205229949
			11'd552: out = 32'b00000000000000001000000000011101; // input=0.53955078125, output=1.00089285236
			11'd553: out = 32'b00000000000000000111111111110111; // input=0.54052734375, output=0.999732543114
			11'd554: out = 32'b00000000000000000111111111010001; // input=0.54150390625, output=0.998571368249
			11'd555: out = 32'b00000000000000000111111110101011; // input=0.54248046875, output=0.99740932426
			11'd556: out = 32'b00000000000000000111111110000101; // input=0.54345703125, output=0.996246407619
			11'd557: out = 32'b00000000000000000111111101011111; // input=0.54443359375, output=0.995082614781
			11'd558: out = 32'b00000000000000000111111100111001; // input=0.54541015625, output=0.993917942183
			11'd559: out = 32'b00000000000000000111111100010011; // input=0.54638671875, output=0.992752386243
			11'd560: out = 32'b00000000000000000111111011101100; // input=0.54736328125, output=0.991585943361
			11'd561: out = 32'b00000000000000000111111011000110; // input=0.54833984375, output=0.990418609919
			11'd562: out = 32'b00000000000000000111111010100000; // input=0.54931640625, output=0.989250382279
			11'd563: out = 32'b00000000000000000111111001111001; // input=0.55029296875, output=0.988081256785
			11'd564: out = 32'b00000000000000000111111001010011; // input=0.55126953125, output=0.986911229762
			11'd565: out = 32'b00000000000000000111111000101101; // input=0.55224609375, output=0.985740297517
			11'd566: out = 32'b00000000000000000111111000000110; // input=0.55322265625, output=0.984568456334
			11'd567: out = 32'b00000000000000000111110111100000; // input=0.55419921875, output=0.983395702482
			11'd568: out = 32'b00000000000000000111110110111001; // input=0.55517578125, output=0.982222032208
			11'd569: out = 32'b00000000000000000111110110010011; // input=0.55615234375, output=0.98104744174
			11'd570: out = 32'b00000000000000000111110101101100; // input=0.55712890625, output=0.979871927286
			11'd571: out = 32'b00000000000000000111110101000110; // input=0.55810546875, output=0.978695485033
			11'd572: out = 32'b00000000000000000111110100011111; // input=0.55908203125, output=0.977518111149
			11'd573: out = 32'b00000000000000000111110011111001; // input=0.56005859375, output=0.976339801781
			11'd574: out = 32'b00000000000000000111110011010010; // input=0.56103515625, output=0.975160553056
			11'd575: out = 32'b00000000000000000111110010101011; // input=0.56201171875, output=0.973980361079
			11'd576: out = 32'b00000000000000000111110010000101; // input=0.56298828125, output=0.972799221937
			11'd577: out = 32'b00000000000000000111110001011110; // input=0.56396484375, output=0.971617131693
			11'd578: out = 32'b00000000000000000111110000110111; // input=0.56494140625, output=0.97043408639
			11'd579: out = 32'b00000000000000000111110000010000; // input=0.56591796875, output=0.96925008205
			11'd580: out = 32'b00000000000000000111101111101010; // input=0.56689453125, output=0.968065114672
			11'd581: out = 32'b00000000000000000111101111000011; // input=0.56787109375, output=0.966879180235
			11'd582: out = 32'b00000000000000000111101110011100; // input=0.56884765625, output=0.965692274695
			11'd583: out = 32'b00000000000000000111101101110101; // input=0.56982421875, output=0.964504393987
			11'd584: out = 32'b00000000000000000111101101001110; // input=0.57080078125, output=0.963315534023
			11'd585: out = 32'b00000000000000000111101100100111; // input=0.57177734375, output=0.962125690692
			11'd586: out = 32'b00000000000000000111101100000000; // input=0.57275390625, output=0.960934859862
			11'd587: out = 32'b00000000000000000111101011011001; // input=0.57373046875, output=0.959743037376
			11'd588: out = 32'b00000000000000000111101010110010; // input=0.57470703125, output=0.958550219057
			11'd589: out = 32'b00000000000000000111101010001011; // input=0.57568359375, output=0.957356400702
			11'd590: out = 32'b00000000000000000111101001100100; // input=0.57666015625, output=0.956161578087
			11'd591: out = 32'b00000000000000000111101000111100; // input=0.57763671875, output=0.954965746961
			11'd592: out = 32'b00000000000000000111101000010101; // input=0.57861328125, output=0.953768903054
			11'd593: out = 32'b00000000000000000111100111101110; // input=0.57958984375, output=0.952571042068
			11'd594: out = 32'b00000000000000000111100111000111; // input=0.58056640625, output=0.951372159683
			11'd595: out = 32'b00000000000000000111100110011111; // input=0.58154296875, output=0.950172251554
			11'd596: out = 32'b00000000000000000111100101111000; // input=0.58251953125, output=0.948971313313
			11'd597: out = 32'b00000000000000000111100101010001; // input=0.58349609375, output=0.947769340563
			11'd598: out = 32'b00000000000000000111100100101001; // input=0.58447265625, output=0.946566328888
			11'd599: out = 32'b00000000000000000111100100000010; // input=0.58544921875, output=0.945362273841
			11'd600: out = 32'b00000000000000000111100011011010; // input=0.58642578125, output=0.944157170955
			11'd601: out = 32'b00000000000000000111100010110011; // input=0.58740234375, output=0.942951015732
			11'd602: out = 32'b00000000000000000111100010001011; // input=0.58837890625, output=0.941743803654
			11'd603: out = 32'b00000000000000000111100001100011; // input=0.58935546875, output=0.940535530172
			11'd604: out = 32'b00000000000000000111100000111100; // input=0.59033203125, output=0.939326190713
			11'd605: out = 32'b00000000000000000111100000010100; // input=0.59130859375, output=0.938115780679
			11'd606: out = 32'b00000000000000000111011111101100; // input=0.59228515625, output=0.936904295441
			11'd607: out = 32'b00000000000000000111011111000101; // input=0.59326171875, output=0.935691730348
			11'd608: out = 32'b00000000000000000111011110011101; // input=0.59423828125, output=0.934478080718
			11'd609: out = 32'b00000000000000000111011101110101; // input=0.59521484375, output=0.933263341845
			11'd610: out = 32'b00000000000000000111011101001101; // input=0.59619140625, output=0.932047508992
			11'd611: out = 32'b00000000000000000111011100100101; // input=0.59716796875, output=0.930830577396
			11'd612: out = 32'b00000000000000000111011011111110; // input=0.59814453125, output=0.929612542267
			11'd613: out = 32'b00000000000000000111011011010110; // input=0.59912109375, output=0.928393398785
			11'd614: out = 32'b00000000000000000111011010101110; // input=0.60009765625, output=0.9271731421
			11'd615: out = 32'b00000000000000000111011010000110; // input=0.60107421875, output=0.925951767338
			11'd616: out = 32'b00000000000000000111011001011110; // input=0.60205078125, output=0.924729269591
			11'd617: out = 32'b00000000000000000111011000110101; // input=0.60302734375, output=0.923505643923
			11'd618: out = 32'b00000000000000000111011000001101; // input=0.60400390625, output=0.922280885371
			11'd619: out = 32'b00000000000000000111010111100101; // input=0.60498046875, output=0.92105498894
			11'd620: out = 32'b00000000000000000111010110111101; // input=0.60595703125, output=0.919827949604
			11'd621: out = 32'b00000000000000000111010110010101; // input=0.60693359375, output=0.918599762308
			11'd622: out = 32'b00000000000000000111010101101100; // input=0.60791015625, output=0.917370421967
			11'd623: out = 32'b00000000000000000111010101000100; // input=0.60888671875, output=0.916139923464
			11'd624: out = 32'b00000000000000000111010100011100; // input=0.60986328125, output=0.91490826165
			11'd625: out = 32'b00000000000000000111010011110011; // input=0.61083984375, output=0.913675431347
			11'd626: out = 32'b00000000000000000111010011001011; // input=0.61181640625, output=0.912441427344
			11'd627: out = 32'b00000000000000000111010010100010; // input=0.61279296875, output=0.911206244396
			11'd628: out = 32'b00000000000000000111010001111010; // input=0.61376953125, output=0.90996987723
			11'd629: out = 32'b00000000000000000111010001010001; // input=0.61474609375, output=0.908732320536
			11'd630: out = 32'b00000000000000000111010000101001; // input=0.61572265625, output=0.907493568975
			11'd631: out = 32'b00000000000000000111010000000000; // input=0.61669921875, output=0.906253617171
			11'd632: out = 32'b00000000000000000111001111010111; // input=0.61767578125, output=0.905012459718
			11'd633: out = 32'b00000000000000000111001110101111; // input=0.61865234375, output=0.903770091174
			11'd634: out = 32'b00000000000000000111001110000110; // input=0.61962890625, output=0.902526506063
			11'd635: out = 32'b00000000000000000111001101011101; // input=0.62060546875, output=0.901281698877
			11'd636: out = 32'b00000000000000000111001100110100; // input=0.62158203125, output=0.90003566407
			11'd637: out = 32'b00000000000000000111001100001011; // input=0.62255859375, output=0.898788396062
			11'd638: out = 32'b00000000000000000111001011100011; // input=0.62353515625, output=0.89753988924
			11'd639: out = 32'b00000000000000000111001010111010; // input=0.62451171875, output=0.896290137952
			11'd640: out = 32'b00000000000000000111001010010001; // input=0.62548828125, output=0.895039136512
			11'd641: out = 32'b00000000000000000111001001101000; // input=0.62646484375, output=0.893786879197
			11'd642: out = 32'b00000000000000000111001000111111; // input=0.62744140625, output=0.892533360247
			11'd643: out = 32'b00000000000000000111001000010101; // input=0.62841796875, output=0.891278573866
			11'd644: out = 32'b00000000000000000111000111101100; // input=0.62939453125, output=0.89002251422
			11'd645: out = 32'b00000000000000000111000111000011; // input=0.63037109375, output=0.888765175437
			11'd646: out = 32'b00000000000000000111000110011010; // input=0.63134765625, output=0.887506551607
			11'd647: out = 32'b00000000000000000111000101110001; // input=0.63232421875, output=0.886246636783
			11'd648: out = 32'b00000000000000000111000101000111; // input=0.63330078125, output=0.884985424977
			11'd649: out = 32'b00000000000000000111000100011110; // input=0.63427734375, output=0.883722910163
			11'd650: out = 32'b00000000000000000111000011110100; // input=0.63525390625, output=0.882459086276
			11'd651: out = 32'b00000000000000000111000011001011; // input=0.63623046875, output=0.881193947211
			11'd652: out = 32'b00000000000000000111000010100001; // input=0.63720703125, output=0.879927486821
			11'd653: out = 32'b00000000000000000111000001111000; // input=0.63818359375, output=0.87865969892
			11'd654: out = 32'b00000000000000000111000001001110; // input=0.63916015625, output=0.877390577281
			11'd655: out = 32'b00000000000000000111000000100101; // input=0.64013671875, output=0.876120115634
			11'd656: out = 32'b00000000000000000110111111111011; // input=0.64111328125, output=0.87484830767
			11'd657: out = 32'b00000000000000000110111111010001; // input=0.64208984375, output=0.873575147036
			11'd658: out = 32'b00000000000000000110111110101000; // input=0.64306640625, output=0.872300627335
			11'd659: out = 32'b00000000000000000110111101111110; // input=0.64404296875, output=0.871024742129
			11'd660: out = 32'b00000000000000000110111101010100; // input=0.64501953125, output=0.869747484936
			11'd661: out = 32'b00000000000000000110111100101010; // input=0.64599609375, output=0.86846884923
			11'd662: out = 32'b00000000000000000110111100000000; // input=0.64697265625, output=0.867188828442
			11'd663: out = 32'b00000000000000000110111011010110; // input=0.64794921875, output=0.865907415954
			11'd664: out = 32'b00000000000000000110111010101100; // input=0.64892578125, output=0.864624605109
			11'd665: out = 32'b00000000000000000110111010000010; // input=0.64990234375, output=0.863340389199
			11'd666: out = 32'b00000000000000000110111001011000; // input=0.65087890625, output=0.862054761472
			11'd667: out = 32'b00000000000000000110111000101110; // input=0.65185546875, output=0.860767715131
			11'd668: out = 32'b00000000000000000110111000000011; // input=0.65283203125, output=0.859479243329
			11'd669: out = 32'b00000000000000000110110111011001; // input=0.65380859375, output=0.858189339174
			11'd670: out = 32'b00000000000000000110110110101111; // input=0.65478515625, output=0.856897995724
			11'd671: out = 32'b00000000000000000110110110000100; // input=0.65576171875, output=0.85560520599
			11'd672: out = 32'b00000000000000000110110101011010; // input=0.65673828125, output=0.854310962935
			11'd673: out = 32'b00000000000000000110110100110000; // input=0.65771484375, output=0.85301525947
			11'd674: out = 32'b00000000000000000110110100000101; // input=0.65869140625, output=0.851718088457
			11'd675: out = 32'b00000000000000000110110011011011; // input=0.65966796875, output=0.850419442709
			11'd676: out = 32'b00000000000000000110110010110000; // input=0.66064453125, output=0.849119314986
			11'd677: out = 32'b00000000000000000110110010000101; // input=0.66162109375, output=0.847817697999
			11'd678: out = 32'b00000000000000000110110001011011; // input=0.66259765625, output=0.846514584405
			11'd679: out = 32'b00000000000000000110110000110000; // input=0.66357421875, output=0.845209966809
			11'd680: out = 32'b00000000000000000110110000000101; // input=0.66455078125, output=0.843903837763
			11'd681: out = 32'b00000000000000000110101111011010; // input=0.66552734375, output=0.842596189766
			11'd682: out = 32'b00000000000000000110101110101111; // input=0.66650390625, output=0.841287015262
			11'd683: out = 32'b00000000000000000110101110000100; // input=0.66748046875, output=0.839976306642
			11'd684: out = 32'b00000000000000000110101101011001; // input=0.66845703125, output=0.838664056239
			11'd685: out = 32'b00000000000000000110101100101110; // input=0.66943359375, output=0.837350256332
			11'd686: out = 32'b00000000000000000110101100000011; // input=0.67041015625, output=0.836034899144
			11'd687: out = 32'b00000000000000000110101011011000; // input=0.67138671875, output=0.83471797684
			11'd688: out = 32'b00000000000000000110101010101101; // input=0.67236328125, output=0.833399481527
			11'd689: out = 32'b00000000000000000110101010000010; // input=0.67333984375, output=0.832079405255
			11'd690: out = 32'b00000000000000000110101001010110; // input=0.67431640625, output=0.830757740015
			11'd691: out = 32'b00000000000000000110101000101011; // input=0.67529296875, output=0.829434477737
			11'd692: out = 32'b00000000000000000110100111111111; // input=0.67626953125, output=0.828109610293
			11'd693: out = 32'b00000000000000000110100111010100; // input=0.67724609375, output=0.826783129494
			11'd694: out = 32'b00000000000000000110100110101001; // input=0.67822265625, output=0.825455027087
			11'd695: out = 32'b00000000000000000110100101111101; // input=0.67919921875, output=0.824125294761
			11'd696: out = 32'b00000000000000000110100101010001; // input=0.68017578125, output=0.82279392414
			11'd697: out = 32'b00000000000000000110100100100110; // input=0.68115234375, output=0.821460906784
			11'd698: out = 32'b00000000000000000110100011111010; // input=0.68212890625, output=0.820126234191
			11'd699: out = 32'b00000000000000000110100011001110; // input=0.68310546875, output=0.818789897792
			11'd700: out = 32'b00000000000000000110100010100010; // input=0.68408203125, output=0.817451888955
			11'd701: out = 32'b00000000000000000110100001110110; // input=0.68505859375, output=0.81611219898
			11'd702: out = 32'b00000000000000000110100001001010; // input=0.68603515625, output=0.814770819101
			11'd703: out = 32'b00000000000000000110100000011110; // input=0.68701171875, output=0.813427740483
			11'd704: out = 32'b00000000000000000110011111110010; // input=0.68798828125, output=0.812082954226
			11'd705: out = 32'b00000000000000000110011111000110; // input=0.68896484375, output=0.810736451356
			11'd706: out = 32'b00000000000000000110011110011010; // input=0.68994140625, output=0.809388222833
			11'd707: out = 32'b00000000000000000110011101101110; // input=0.69091796875, output=0.808038259545
			11'd708: out = 32'b00000000000000000110011101000010; // input=0.69189453125, output=0.806686552309
			11'd709: out = 32'b00000000000000000110011100010101; // input=0.69287109375, output=0.805333091869
			11'd710: out = 32'b00000000000000000110011011101001; // input=0.69384765625, output=0.803977868896
			11'd711: out = 32'b00000000000000000110011010111100; // input=0.69482421875, output=0.802620873988
			11'd712: out = 32'b00000000000000000110011010010000; // input=0.69580078125, output=0.801262097667
			11'd713: out = 32'b00000000000000000110011001100011; // input=0.69677734375, output=0.799901530381
			11'd714: out = 32'b00000000000000000110011000110111; // input=0.69775390625, output=0.798539162501
			11'd715: out = 32'b00000000000000000110011000001010; // input=0.69873046875, output=0.79717498432
			11'd716: out = 32'b00000000000000000110010111011101; // input=0.69970703125, output=0.795808986053
			11'd717: out = 32'b00000000000000000110010110110000; // input=0.70068359375, output=0.794441157837
			11'd718: out = 32'b00000000000000000110010110000011; // input=0.70166015625, output=0.793071489728
			11'd719: out = 32'b00000000000000000110010101010110; // input=0.70263671875, output=0.791699971702
			11'd720: out = 32'b00000000000000000110010100101001; // input=0.70361328125, output=0.790326593651
			11'd721: out = 32'b00000000000000000110010011111100; // input=0.70458984375, output=0.788951345388
			11'd722: out = 32'b00000000000000000110010011001111; // input=0.70556640625, output=0.787574216638
			11'd723: out = 32'b00000000000000000110010010100010; // input=0.70654296875, output=0.786195197045
			11'd724: out = 32'b00000000000000000110010001110101; // input=0.70751953125, output=0.784814276165
			11'd725: out = 32'b00000000000000000110010001000111; // input=0.70849609375, output=0.783431443467
			11'd726: out = 32'b00000000000000000110010000011010; // input=0.70947265625, output=0.782046688334
			11'd727: out = 32'b00000000000000000110001111101101; // input=0.71044921875, output=0.78066000006
			11'd728: out = 32'b00000000000000000110001110111111; // input=0.71142578125, output=0.779271367848
			11'd729: out = 32'b00000000000000000110001110010010; // input=0.71240234375, output=0.77788078081
			11'd730: out = 32'b00000000000000000110001101100100; // input=0.71337890625, output=0.776488227967
			11'd731: out = 32'b00000000000000000110001100110110; // input=0.71435546875, output=0.775093698247
			11'd732: out = 32'b00000000000000000110001100001001; // input=0.71533203125, output=0.773697180483
			11'd733: out = 32'b00000000000000000110001011011011; // input=0.71630859375, output=0.772298663413
			11'd734: out = 32'b00000000000000000110001010101101; // input=0.71728515625, output=0.770898135678
			11'd735: out = 32'b00000000000000000110001001111111; // input=0.71826171875, output=0.769495585822
			11'd736: out = 32'b00000000000000000110001001010001; // input=0.71923828125, output=0.768091002289
			11'd737: out = 32'b00000000000000000110001000100011; // input=0.72021484375, output=0.766684373425
			11'd738: out = 32'b00000000000000000110000111110101; // input=0.72119140625, output=0.765275687473
			11'd739: out = 32'b00000000000000000110000111000110; // input=0.72216796875, output=0.763864932573
			11'd740: out = 32'b00000000000000000110000110011000; // input=0.72314453125, output=0.762452096763
			11'd741: out = 32'b00000000000000000110000101101010; // input=0.72412109375, output=0.761037167974
			11'd742: out = 32'b00000000000000000110000100111011; // input=0.72509765625, output=0.759620134032
			11'd743: out = 32'b00000000000000000110000100001101; // input=0.72607421875, output=0.758200982654
			11'd744: out = 32'b00000000000000000110000011011110; // input=0.72705078125, output=0.756779701448
			11'd745: out = 32'b00000000000000000110000010110000; // input=0.72802734375, output=0.755356277913
			11'd746: out = 32'b00000000000000000110000010000001; // input=0.72900390625, output=0.753930699434
			11'd747: out = 32'b00000000000000000110000001010010; // input=0.72998046875, output=0.752502953285
			11'd748: out = 32'b00000000000000000110000000100011; // input=0.73095703125, output=0.751073026622
			11'd749: out = 32'b00000000000000000101111111110100; // input=0.73193359375, output=0.749640906488
			11'd750: out = 32'b00000000000000000101111111000101; // input=0.73291015625, output=0.748206579806
			11'd751: out = 32'b00000000000000000101111110010110; // input=0.73388671875, output=0.746770033382
			11'd752: out = 32'b00000000000000000101111101100111; // input=0.73486328125, output=0.745331253898
			11'd753: out = 32'b00000000000000000101111100111000; // input=0.73583984375, output=0.743890227917
			11'd754: out = 32'b00000000000000000101111100001001; // input=0.73681640625, output=0.742446941877
			11'd755: out = 32'b00000000000000000101111011011001; // input=0.73779296875, output=0.741001382088
			11'd756: out = 32'b00000000000000000101111010101010; // input=0.73876953125, output=0.739553534736
			11'd757: out = 32'b00000000000000000101111001111010; // input=0.73974609375, output=0.738103385877
			11'd758: out = 32'b00000000000000000101111001001011; // input=0.74072265625, output=0.736650921436
			11'd759: out = 32'b00000000000000000101111000011011; // input=0.74169921875, output=0.735196127207
			11'd760: out = 32'b00000000000000000101110111101011; // input=0.74267578125, output=0.733738988847
			11'd761: out = 32'b00000000000000000101110110111011; // input=0.74365234375, output=0.73227949188
			11'd762: out = 32'b00000000000000000101110110001011; // input=0.74462890625, output=0.730817621692
			11'd763: out = 32'b00000000000000000101110101011011; // input=0.74560546875, output=0.729353363528
			11'd764: out = 32'b00000000000000000101110100101011; // input=0.74658203125, output=0.727886702492
			11'd765: out = 32'b00000000000000000101110011111011; // input=0.74755859375, output=0.726417623546
			11'd766: out = 32'b00000000000000000101110011001011; // input=0.74853515625, output=0.724946111505
			11'd767: out = 32'b00000000000000000101110010011011; // input=0.74951171875, output=0.723472151039
			11'd768: out = 32'b00000000000000000101110001101010; // input=0.75048828125, output=0.721995726665
			11'd769: out = 32'b00000000000000000101110000111010; // input=0.75146484375, output=0.720516822751
			11'd770: out = 32'b00000000000000000101110000001001; // input=0.75244140625, output=0.719035423513
			11'd771: out = 32'b00000000000000000101101111011001; // input=0.75341796875, output=0.717551513008
			11'd772: out = 32'b00000000000000000101101110101000; // input=0.75439453125, output=0.716065075138
			11'd773: out = 32'b00000000000000000101101101110111; // input=0.75537109375, output=0.714576093643
			11'd774: out = 32'b00000000000000000101101101000110; // input=0.75634765625, output=0.713084552103
			11'd775: out = 32'b00000000000000000101101100010101; // input=0.75732421875, output=0.711590433931
			11'd776: out = 32'b00000000000000000101101011100100; // input=0.75830078125, output=0.710093722376
			11'd777: out = 32'b00000000000000000101101010110011; // input=0.75927734375, output=0.708594400515
			11'd778: out = 32'b00000000000000000101101010000010; // input=0.76025390625, output=0.707092451256
			11'd779: out = 32'b00000000000000000101101001010001; // input=0.76123046875, output=0.70558785733
			11'd780: out = 32'b00000000000000000101101000011111; // input=0.76220703125, output=0.704080601293
			11'd781: out = 32'b00000000000000000101100111101110; // input=0.76318359375, output=0.702570665524
			11'd782: out = 32'b00000000000000000101100110111100; // input=0.76416015625, output=0.701058032216
			11'd783: out = 32'b00000000000000000101100110001011; // input=0.76513671875, output=0.699542683381
			11'd784: out = 32'b00000000000000000101100101011001; // input=0.76611328125, output=0.698024600842
			11'd785: out = 32'b00000000000000000101100100100111; // input=0.76708984375, output=0.696503766233
			11'd786: out = 32'b00000000000000000101100011110101; // input=0.76806640625, output=0.694980160996
			11'd787: out = 32'b00000000000000000101100011000011; // input=0.76904296875, output=0.693453766377
			11'd788: out = 32'b00000000000000000101100010010001; // input=0.77001953125, output=0.691924563422
			11'd789: out = 32'b00000000000000000101100001011111; // input=0.77099609375, output=0.690392532978
			11'd790: out = 32'b00000000000000000101100000101100; // input=0.77197265625, output=0.688857655687
			11'd791: out = 32'b00000000000000000101011111111010; // input=0.77294921875, output=0.687319911983
			11'd792: out = 32'b00000000000000000101011111001000; // input=0.77392578125, output=0.685779282091
			11'd793: out = 32'b00000000000000000101011110010101; // input=0.77490234375, output=0.684235746018
			11'd794: out = 32'b00000000000000000101011101100010; // input=0.77587890625, output=0.68268928356
			11'd795: out = 32'b00000000000000000101011100110000; // input=0.77685546875, output=0.681139874289
			11'd796: out = 32'b00000000000000000101011011111101; // input=0.77783203125, output=0.679587497552
			11'd797: out = 32'b00000000000000000101011011001010; // input=0.77880859375, output=0.678032132473
			11'd798: out = 32'b00000000000000000101011010010111; // input=0.77978515625, output=0.676473757941
			11'd799: out = 32'b00000000000000000101011001100100; // input=0.78076171875, output=0.674912352614
			11'd800: out = 32'b00000000000000000101011000110000; // input=0.78173828125, output=0.67334789491
			11'd801: out = 32'b00000000000000000101010111111101; // input=0.78271484375, output=0.671780363006
			11'd802: out = 32'b00000000000000000101010111001001; // input=0.78369140625, output=0.670209734833
			11'd803: out = 32'b00000000000000000101010110010110; // input=0.78466796875, output=0.668635988073
			11'd804: out = 32'b00000000000000000101010101100010; // input=0.78564453125, output=0.667059100154
			11'd805: out = 32'b00000000000000000101010100101110; // input=0.78662109375, output=0.665479048247
			11'd806: out = 32'b00000000000000000101010011111011; // input=0.78759765625, output=0.663895809262
			11'd807: out = 32'b00000000000000000101010011000111; // input=0.78857421875, output=0.662309359842
			11'd808: out = 32'b00000000000000000101010010010010; // input=0.78955078125, output=0.660719676359
			11'd809: out = 32'b00000000000000000101010001011110; // input=0.79052734375, output=0.659126734912
			11'd810: out = 32'b00000000000000000101010000101010; // input=0.79150390625, output=0.657530511322
			11'd811: out = 32'b00000000000000000101001111110110; // input=0.79248046875, output=0.655930981122
			11'd812: out = 32'b00000000000000000101001111000001; // input=0.79345703125, output=0.654328119562
			11'd813: out = 32'b00000000000000000101001110001100; // input=0.79443359375, output=0.652721901594
			11'd814: out = 32'b00000000000000000101001101011000; // input=0.79541015625, output=0.651112301876
			11'd815: out = 32'b00000000000000000101001100100011; // input=0.79638671875, output=0.649499294759
			11'd816: out = 32'b00000000000000000101001011101110; // input=0.79736328125, output=0.647882854289
			11'd817: out = 32'b00000000000000000101001010111001; // input=0.79833984375, output=0.646262954198
			11'd818: out = 32'b00000000000000000101001010000100; // input=0.79931640625, output=0.644639567897
			11'd819: out = 32'b00000000000000000101001001001110; // input=0.80029296875, output=0.643012668475
			11'd820: out = 32'b00000000000000000101001000011001; // input=0.80126953125, output=0.64138222869
			11'd821: out = 32'b00000000000000000101000111100011; // input=0.80224609375, output=0.639748220967
			11'd822: out = 32'b00000000000000000101000110101110; // input=0.80322265625, output=0.638110617386
			11'd823: out = 32'b00000000000000000101000101111000; // input=0.80419921875, output=0.636469389683
			11'd824: out = 32'b00000000000000000101000101000010; // input=0.80517578125, output=0.634824509238
			11'd825: out = 32'b00000000000000000101000100001100; // input=0.80615234375, output=0.633175947074
			11'd826: out = 32'b00000000000000000101000011010110; // input=0.80712890625, output=0.631523673845
			11'd827: out = 32'b00000000000000000101000010100000; // input=0.80810546875, output=0.629867659836
			11'd828: out = 32'b00000000000000000101000001101001; // input=0.80908203125, output=0.62820787495
			11'd829: out = 32'b00000000000000000101000000110011; // input=0.81005859375, output=0.626544288707
			11'd830: out = 32'b00000000000000000100111111111100; // input=0.81103515625, output=0.62487687023
			11'd831: out = 32'b00000000000000000100111111000101; // input=0.81201171875, output=0.623205588247
			11'd832: out = 32'b00000000000000000100111110001110; // input=0.81298828125, output=0.621530411074
			11'd833: out = 32'b00000000000000000100111101010111; // input=0.81396484375, output=0.619851306615
			11'd834: out = 32'b00000000000000000100111100100000; // input=0.81494140625, output=0.61816824235
			11'd835: out = 32'b00000000000000000100111011101001; // input=0.81591796875, output=0.616481185331
			11'd836: out = 32'b00000000000000000100111010110001; // input=0.81689453125, output=0.614790102169
			11'd837: out = 32'b00000000000000000100111001111010; // input=0.81787109375, output=0.61309495903
			11'd838: out = 32'b00000000000000000100111001000010; // input=0.81884765625, output=0.611395721625
			11'd839: out = 32'b00000000000000000100111000001010; // input=0.81982421875, output=0.6096923552
			11'd840: out = 32'b00000000000000000100110111010010; // input=0.82080078125, output=0.607984824531
			11'd841: out = 32'b00000000000000000100110110011010; // input=0.82177734375, output=0.60627309391
			11'd842: out = 32'b00000000000000000100110101100010; // input=0.82275390625, output=0.60455712714
			11'd843: out = 32'b00000000000000000100110100101010; // input=0.82373046875, output=0.602836887524
			11'd844: out = 32'b00000000000000000100110011110001; // input=0.82470703125, output=0.601112337854
			11'd845: out = 32'b00000000000000000100110010111001; // input=0.82568359375, output=0.599383440402
			11'd846: out = 32'b00000000000000000100110010000000; // input=0.82666015625, output=0.597650156911
			11'd847: out = 32'b00000000000000000100110001000111; // input=0.82763671875, output=0.595912448581
			11'd848: out = 32'b00000000000000000100110000001110; // input=0.82861328125, output=0.594170276064
			11'd849: out = 32'b00000000000000000100101111010101; // input=0.82958984375, output=0.592423599447
			11'd850: out = 32'b00000000000000000100101110011011; // input=0.83056640625, output=0.590672378243
			11'd851: out = 32'b00000000000000000100101101100010; // input=0.83154296875, output=0.588916571382
			11'd852: out = 32'b00000000000000000100101100101000; // input=0.83251953125, output=0.587156137194
			11'd853: out = 32'b00000000000000000100101011101110; // input=0.83349609375, output=0.585391033401
			11'd854: out = 32'b00000000000000000100101010110100; // input=0.83447265625, output=0.583621217101
			11'd855: out = 32'b00000000000000000100101001111010; // input=0.83544921875, output=0.58184664476
			11'd856: out = 32'b00000000000000000100101001000000; // input=0.83642578125, output=0.580067272194
			11'd857: out = 32'b00000000000000000100101000000101; // input=0.83740234375, output=0.578283054556
			11'd858: out = 32'b00000000000000000100100111001011; // input=0.83837890625, output=0.576493946324
			11'd859: out = 32'b00000000000000000100100110010000; // input=0.83935546875, output=0.574699901288
			11'd860: out = 32'b00000000000000000100100101010101; // input=0.84033203125, output=0.572900872529
			11'd861: out = 32'b00000000000000000100100100011010; // input=0.84130859375, output=0.571096812411
			11'd862: out = 32'b00000000000000000100100011011110; // input=0.84228515625, output=0.569287672562
			11'd863: out = 32'b00000000000000000100100010100011; // input=0.84326171875, output=0.567473403856
			11'd864: out = 32'b00000000000000000100100001100111; // input=0.84423828125, output=0.565653956402
			11'd865: out = 32'b00000000000000000100100000101100; // input=0.84521484375, output=0.563829279521
			11'd866: out = 32'b00000000000000000100011111110000; // input=0.84619140625, output=0.561999321734
			11'd867: out = 32'b00000000000000000100011110110011; // input=0.84716796875, output=0.560164030741
			11'd868: out = 32'b00000000000000000100011101110111; // input=0.84814453125, output=0.558323353402
			11'd869: out = 32'b00000000000000000100011100111011; // input=0.84912109375, output=0.556477235721
			11'd870: out = 32'b00000000000000000100011011111110; // input=0.85009765625, output=0.554625622823
			11'd871: out = 32'b00000000000000000100011011000001; // input=0.85107421875, output=0.552768458938
			11'd872: out = 32'b00000000000000000100011010000100; // input=0.85205078125, output=0.550905687375
			11'd873: out = 32'b00000000000000000100011001000111; // input=0.85302734375, output=0.549037250506
			11'd874: out = 32'b00000000000000000100011000001001; // input=0.85400390625, output=0.547163089742
			11'd875: out = 32'b00000000000000000100010111001100; // input=0.85498046875, output=0.545283145509
			11'd876: out = 32'b00000000000000000100010110001110; // input=0.85595703125, output=0.543397357226
			11'd877: out = 32'b00000000000000000100010101010000; // input=0.85693359375, output=0.541505663281
			11'd878: out = 32'b00000000000000000100010100010010; // input=0.85791015625, output=0.539608001008
			11'd879: out = 32'b00000000000000000100010011010011; // input=0.85888671875, output=0.537704306657
			11'd880: out = 32'b00000000000000000100010010010101; // input=0.85986328125, output=0.535794515372
			11'd881: out = 32'b00000000000000000100010001010110; // input=0.86083984375, output=0.533878561162
			11'd882: out = 32'b00000000000000000100010000010111; // input=0.86181640625, output=0.531956376874
			11'd883: out = 32'b00000000000000000100001111011000; // input=0.86279296875, output=0.530027894162
			11'd884: out = 32'b00000000000000000100001110011001; // input=0.86376953125, output=0.528093043461
			11'd885: out = 32'b00000000000000000100001101011001; // input=0.86474609375, output=0.526151753951
			11'd886: out = 32'b00000000000000000100001100011001; // input=0.86572265625, output=0.524203953531
			11'd887: out = 32'b00000000000000000100001011011001; // input=0.86669921875, output=0.522249568781
			11'd888: out = 32'b00000000000000000100001010011001; // input=0.86767578125, output=0.520288524932
			11'd889: out = 32'b00000000000000000100001001011000; // input=0.86865234375, output=0.51832074583
			11'd890: out = 32'b00000000000000000100001000011000; // input=0.86962890625, output=0.516346153897
			11'd891: out = 32'b00000000000000000100000111010111; // input=0.87060546875, output=0.514364670098
			11'd892: out = 32'b00000000000000000100000110010110; // input=0.87158203125, output=0.5123762139
			11'd893: out = 32'b00000000000000000100000101010100; // input=0.87255859375, output=0.51038070323
			11'd894: out = 32'b00000000000000000100000100010011; // input=0.87353515625, output=0.508378054438
			11'd895: out = 32'b00000000000000000100000011010001; // input=0.87451171875, output=0.506368182252
			11'd896: out = 32'b00000000000000000100000010001111; // input=0.87548828125, output=0.504350999733
			11'd897: out = 32'b00000000000000000100000001001100; // input=0.87646484375, output=0.502326418228
			11'd898: out = 32'b00000000000000000100000000001010; // input=0.87744140625, output=0.500294347326
			11'd899: out = 32'b00000000000000000011111111000111; // input=0.87841796875, output=0.498254694808
			11'd900: out = 32'b00000000000000000011111110000100; // input=0.87939453125, output=0.496207366591
			11'd901: out = 32'b00000000000000000011111101000000; // input=0.88037109375, output=0.494152266683
			11'd902: out = 32'b00000000000000000011111011111101; // input=0.88134765625, output=0.492089297121
			11'd903: out = 32'b00000000000000000011111010111001; // input=0.88232421875, output=0.490018357918
			11'd904: out = 32'b00000000000000000011111001110101; // input=0.88330078125, output=0.487939347004
			11'd905: out = 32'b00000000000000000011111000110000; // input=0.88427734375, output=0.485852160163
			11'd906: out = 32'b00000000000000000011110111101100; // input=0.88525390625, output=0.483756690969
			11'd907: out = 32'b00000000000000000011110110100111; // input=0.88623046875, output=0.481652830723
			11'd908: out = 32'b00000000000000000011110101100010; // input=0.88720703125, output=0.479540468383
			11'd909: out = 32'b00000000000000000011110100011100; // input=0.88818359375, output=0.47741949049
			11'd910: out = 32'b00000000000000000011110011010110; // input=0.88916015625, output=0.475289781097
			11'd911: out = 32'b00000000000000000011110010010000; // input=0.89013671875, output=0.473151221691
			11'd912: out = 32'b00000000000000000011110001001010; // input=0.89111328125, output=0.471003691115
			11'd913: out = 32'b00000000000000000011110000000011; // input=0.89208984375, output=0.468847065479
			11'd914: out = 32'b00000000000000000011101110111100; // input=0.89306640625, output=0.46668121808
			11'd915: out = 32'b00000000000000000011101101110101; // input=0.89404296875, output=0.464506019307
			11'd916: out = 32'b00000000000000000011101100101101; // input=0.89501953125, output=0.462321336549
			11'd917: out = 32'b00000000000000000011101011100101; // input=0.89599609375, output=0.460127034094
			11'd918: out = 32'b00000000000000000011101010011101; // input=0.89697265625, output=0.457922973032
			11'd919: out = 32'b00000000000000000011101001010101; // input=0.89794921875, output=0.455709011145
			11'd920: out = 32'b00000000000000000011101000001100; // input=0.89892578125, output=0.453485002794
			11'd921: out = 32'b00000000000000000011100111000011; // input=0.89990234375, output=0.451250798807
			11'd922: out = 32'b00000000000000000011100101111001; // input=0.90087890625, output=0.449006246355
			11'd923: out = 32'b00000000000000000011100100101111; // input=0.90185546875, output=0.446751188828
			11'd924: out = 32'b00000000000000000011100011100101; // input=0.90283203125, output=0.444485465699
			11'd925: out = 32'b00000000000000000011100010011010; // input=0.90380859375, output=0.442208912389
			11'd926: out = 32'b00000000000000000011100001001111; // input=0.90478515625, output=0.439921360122
			11'd927: out = 32'b00000000000000000011100000000100; // input=0.90576171875, output=0.437622635771
			11'd928: out = 32'b00000000000000000011011110111000; // input=0.90673828125, output=0.435312561704
			11'd929: out = 32'b00000000000000000011011101101100; // input=0.90771484375, output=0.432990955614
			11'd930: out = 32'b00000000000000000011011100100000; // input=0.90869140625, output=0.430657630348
			11'd931: out = 32'b00000000000000000011011011010011; // input=0.90966796875, output=0.428312393723
			11'd932: out = 32'b00000000000000000011011010000110; // input=0.91064453125, output=0.425955048337
			11'd933: out = 32'b00000000000000000011011000111000; // input=0.91162109375, output=0.423585391365
			11'd934: out = 32'b00000000000000000011010111101010; // input=0.91259765625, output=0.421203214354
			11'd935: out = 32'b00000000000000000011010110011100; // input=0.91357421875, output=0.418808302995
			11'd936: out = 32'b00000000000000000011010101001101; // input=0.91455078125, output=0.416400436898
			11'd937: out = 32'b00000000000000000011010011111101; // input=0.91552734375, output=0.413979389341
			11'd938: out = 32'b00000000000000000011010010101110; // input=0.91650390625, output=0.411544927017
			11'd939: out = 32'b00000000000000000011010001011101; // input=0.91748046875, output=0.409096809761
			11'd940: out = 32'b00000000000000000011010000001101; // input=0.91845703125, output=0.406634790267
			11'd941: out = 32'b00000000000000000011001110111011; // input=0.91943359375, output=0.404158613784
			11'd942: out = 32'b00000000000000000011001101101010; // input=0.92041015625, output=0.401668017804
			11'd943: out = 32'b00000000000000000011001100011000; // input=0.92138671875, output=0.399162731721
			11'd944: out = 32'b00000000000000000011001011000101; // input=0.92236328125, output=0.396642476482
			11'd945: out = 32'b00000000000000000011001001110010; // input=0.92333984375, output=0.394106964214
			11'd946: out = 32'b00000000000000000011001000011111; // input=0.92431640625, output=0.391555897824
			11'd947: out = 32'b00000000000000000011000111001010; // input=0.92529296875, output=0.388988970587
			11'd948: out = 32'b00000000000000000011000101110110; // input=0.92626953125, output=0.386405865698
			11'd949: out = 32'b00000000000000000011000100100001; // input=0.92724609375, output=0.383806255807
			11'd950: out = 32'b00000000000000000011000011001011; // input=0.92822265625, output=0.381189802517
			11'd951: out = 32'b00000000000000000011000001110101; // input=0.92919921875, output=0.378556155859
			11'd952: out = 32'b00000000000000000011000000011110; // input=0.93017578125, output=0.375904953732
			11'd953: out = 32'b00000000000000000010111111000110; // input=0.93115234375, output=0.3732358213
			11'd954: out = 32'b00000000000000000010111101101110; // input=0.93212890625, output=0.370548370363
			11'd955: out = 32'b00000000000000000010111100010101; // input=0.93310546875, output=0.36784219868
			11'd956: out = 32'b00000000000000000010111010111100; // input=0.93408203125, output=0.365116889244
			11'd957: out = 32'b00000000000000000010111001100010; // input=0.93505859375, output=0.362372009518
			11'd958: out = 32'b00000000000000000010111000001000; // input=0.93603515625, output=0.359607110609
			11'd959: out = 32'b00000000000000000010110110101100; // input=0.93701171875, output=0.356821726393
			11'd960: out = 32'b00000000000000000010110101010000; // input=0.93798828125, output=0.354015372576
			11'd961: out = 32'b00000000000000000010110011110100; // input=0.93896484375, output=0.351187545683
			11'd962: out = 32'b00000000000000000010110010010110; // input=0.93994140625, output=0.348337721984
			11'd963: out = 32'b00000000000000000010110000111000; // input=0.94091796875, output=0.345465356329
			11'd964: out = 32'b00000000000000000010101111011001; // input=0.94189453125, output=0.34256988091
			11'd965: out = 32'b00000000000000000010101101111010; // input=0.94287109375, output=0.339650703915
			11'd966: out = 32'b00000000000000000010101100011001; // input=0.94384765625, output=0.336707208087
			11'd967: out = 32'b00000000000000000010101010111000; // input=0.94482421875, output=0.333738749167
			11'd968: out = 32'b00000000000000000010101001010110; // input=0.94580078125, output=0.330744654211
			11'd969: out = 32'b00000000000000000010100111110011; // input=0.94677734375, output=0.327724219773
			11'd970: out = 32'b00000000000000000010100110001111; // input=0.94775390625, output=0.324676709931
			11'd971: out = 32'b00000000000000000010100100101010; // input=0.94873046875, output=0.321601354156
			11'd972: out = 32'b00000000000000000010100011000101; // input=0.94970703125, output=0.318497344988
			11'd973: out = 32'b00000000000000000010100001011110; // input=0.95068359375, output=0.315363835514
			11'd974: out = 32'b00000000000000000010011111110110; // input=0.95166015625, output=0.312199936613
			11'd975: out = 32'b00000000000000000010011110001101; // input=0.95263671875, output=0.309004713959
			11'd976: out = 32'b00000000000000000010011100100100; // input=0.95361328125, output=0.305777184735
			11'd977: out = 32'b00000000000000000010011010111001; // input=0.95458984375, output=0.302516314039
			11'd978: out = 32'b00000000000000000010011001001101; // input=0.95556640625, output=0.299221010939
			11'd979: out = 32'b00000000000000000010010111100000; // input=0.95654296875, output=0.295890124136
			11'd980: out = 32'b00000000000000000010010101110001; // input=0.95751953125, output=0.292522437183
			11'd981: out = 32'b00000000000000000010010100000010; // input=0.95849609375, output=0.289116663208
			11'd982: out = 32'b00000000000000000010010010010001; // input=0.95947265625, output=0.285671439076
			11'd983: out = 32'b00000000000000000010010000011111; // input=0.96044921875, output=0.282185318912
			11'd984: out = 32'b00000000000000000010001110101011; // input=0.96142578125, output=0.278656766898
			11'd985: out = 32'b00000000000000000010001100110110; // input=0.96240234375, output=0.275084149249
			11'd986: out = 32'b00000000000000000010001010111111; // input=0.96337890625, output=0.271465725233
			11'd987: out = 32'b00000000000000000010001001000111; // input=0.96435546875, output=0.267799637122
			11'd988: out = 32'b00000000000000000010000111001110; // input=0.96533203125, output=0.264083898876
			11'd989: out = 32'b00000000000000000010000101010010; // input=0.96630859375, output=0.260316383399
			11'd990: out = 32'b00000000000000000010000011010101; // input=0.96728515625, output=0.256494808104
			11'd991: out = 32'b00000000000000000010000001010110; // input=0.96826171875, output=0.252616718532
			11'd992: out = 32'b00000000000000000001111111010101; // input=0.96923828125, output=0.248679469682
			11'd993: out = 32'b00000000000000000001111101010010; // input=0.97021484375, output=0.244680204644
			11'd994: out = 32'b00000000000000000001111011001100; // input=0.97119140625, output=0.240615830061
			11'd995: out = 32'b00000000000000000001111001000101; // input=0.97216796875, output=0.236482987801
			11'd996: out = 32'b00000000000000000001110110111011; // input=0.97314453125, output=0.232278022117
			11'd997: out = 32'b00000000000000000001110100101111; // input=0.97412109375, output=0.227996941384
			11'd998: out = 32'b00000000000000000001110010100000; // input=0.97509765625, output=0.223635373253
			11'd999: out = 32'b00000000000000000001110000001110; // input=0.97607421875, output=0.219188511821
			11'd1000: out = 32'b00000000000000000001101101111010; // input=0.97705078125, output=0.214651054972
			11'd1001: out = 32'b00000000000000000001101011100010; // input=0.97802734375, output=0.210017129581
			11'd1002: out = 32'b00000000000000000001101001000111; // input=0.97900390625, output=0.20528020156
			11'd1003: out = 32'b00000000000000000001100110101000; // input=0.97998046875, output=0.200432966839
			11'd1004: out = 32'b00000000000000000001100100000101; // input=0.98095703125, output=0.195467218063
			11'd1005: out = 32'b00000000000000000001100001011110; // input=0.98193359375, output=0.19037368008
			11'd1006: out = 32'b00000000000000000001011110110011; // input=0.98291015625, output=0.185141804779
			11'd1007: out = 32'b00000000000000000001011100000010; // input=0.98388671875, output=0.179759512289
			11'd1008: out = 32'b00000000000000000001011001001101; // input=0.98486328125, output=0.17421286033
			11'd1009: out = 32'b00000000000000000001010110010001; // input=0.98583984375, output=0.168485615729
			11'd1010: out = 32'b00000000000000000001010011001111; // input=0.98681640625, output=0.162558690208
			11'd1011: out = 32'b00000000000000000001010000000101; // input=0.98779296875, output=0.15640938387
			11'd1012: out = 32'b00000000000000000001001100110100; // input=0.98876953125, output=0.150010349655
			11'd1013: out = 32'b00000000000000000001001001011001; // input=0.98974609375, output=0.143328141623
			11'd1014: out = 32'b00000000000000000001000101110011; // input=0.99072265625, output=0.136321122325
			11'd1015: out = 32'b00000000000000000001000010000001; // input=0.99169921875, output=0.128936345273
			11'd1016: out = 32'b00000000000000000000111110000000; // input=0.99267578125, output=0.121104722866
			11'd1017: out = 32'b00000000000000000000111001101110; // input=0.99365234375, output=0.112733163685
			11'd1018: out = 32'b00000000000000000000110101000110; // input=0.99462890625, output=0.103690971223
			11'd1019: out = 32'b00000000000000000000110000000001; // input=0.99560546875, output=0.0937843662666
			11'd1020: out = 32'b00000000000000000000101010010110; // input=0.99658203125, output=0.0827032963273
			11'd1021: out = 32'b00000000000000000000100011110010; // input=0.99755859375, output=0.0698913486493
			11'd1022: out = 32'b00000000000000000000011011101110; // input=0.99853515625, output=0.0541331971646
			11'd1023: out = 32'b00000000000000000000010000000000; // input=0.99951171875, output=0.0312512717055
			11'd1024: out = 32'b00000000000000001100100100100000; // input=-0.00048828125, output=1.57128460806
			11'd1025: out = 32'b00000000000000001100100101000000; // input=-0.00146484375, output=1.57226117107
			11'd1026: out = 32'b00000000000000001100100101100000; // input=-0.00244140625, output=1.57323773547
			11'd1027: out = 32'b00000000000000001100100110000000; // input=-0.00341796875, output=1.5742143022
			11'd1028: out = 32'b00000000000000001100100110100000; // input=-0.00439453125, output=1.57519087219
			11'd1029: out = 32'b00000000000000001100100111000000; // input=-0.00537109375, output=1.57616744637
			11'd1030: out = 32'b00000000000000001100100111100000; // input=-0.00634765625, output=1.57714402567
			11'd1031: out = 32'b00000000000000001100101000000000; // input=-0.00732421875, output=1.57812061103
			11'd1032: out = 32'b00000000000000001100101000100000; // input=-0.00830078125, output=1.57909720337
			11'd1033: out = 32'b00000000000000001100101001000000; // input=-0.00927734375, output=1.58007380363
			11'd1034: out = 32'b00000000000000001100101001100000; // input=-0.01025390625, output=1.58105041274
			11'd1035: out = 32'b00000000000000001100101010000000; // input=-0.01123046875, output=1.58202703163
			11'd1036: out = 32'b00000000000000001100101010100000; // input=-0.01220703125, output=1.58300366123
			11'd1037: out = 32'b00000000000000001100101011000000; // input=-0.01318359375, output=1.58398030248
			11'd1038: out = 32'b00000000000000001100101011100000; // input=-0.01416015625, output=1.5849569563
			11'd1039: out = 32'b00000000000000001100101100000000; // input=-0.01513671875, output=1.58593362363
			11'd1040: out = 32'b00000000000000001100101100100000; // input=-0.01611328125, output=1.5869103054
			11'd1041: out = 32'b00000000000000001100101101000000; // input=-0.01708984375, output=1.58788700254
			11'd1042: out = 32'b00000000000000001100101101100000; // input=-0.01806640625, output=1.58886371599
			11'd1043: out = 32'b00000000000000001100101110000000; // input=-0.01904296875, output=1.58984044667
			11'd1044: out = 32'b00000000000000001100101110100000; // input=-0.02001953125, output=1.59081719553
			11'd1045: out = 32'b00000000000000001100101111000000; // input=-0.02099609375, output=1.59179396349
			11'd1046: out = 32'b00000000000000001100101111100000; // input=-0.02197265625, output=1.59277075149
			11'd1047: out = 32'b00000000000000001100110000000000; // input=-0.02294921875, output=1.59374756045
			11'd1048: out = 32'b00000000000000001100110000100000; // input=-0.02392578125, output=1.59472439132
			11'd1049: out = 32'b00000000000000001100110001000000; // input=-0.02490234375, output=1.59570124503
			11'd1050: out = 32'b00000000000000001100110001100000; // input=-0.02587890625, output=1.59667812251
			11'd1051: out = 32'b00000000000000001100110010000000; // input=-0.02685546875, output=1.59765502469
			11'd1052: out = 32'b00000000000000001100110010100000; // input=-0.02783203125, output=1.59863195252
			11'd1053: out = 32'b00000000000000001100110011000000; // input=-0.02880859375, output=1.59960890691
			11'd1054: out = 32'b00000000000000001100110011100000; // input=-0.02978515625, output=1.60058588882
			11'd1055: out = 32'b00000000000000001100110100000000; // input=-0.03076171875, output=1.60156289916
			11'd1056: out = 32'b00000000000000001100110100100000; // input=-0.03173828125, output=1.60253993889
			11'd1057: out = 32'b00000000000000001100110101000000; // input=-0.03271484375, output=1.60351700893
			11'd1058: out = 32'b00000000000000001100110101100000; // input=-0.03369140625, output=1.60449411022
			11'd1059: out = 32'b00000000000000001100110110000000; // input=-0.03466796875, output=1.60547124369
			11'd1060: out = 32'b00000000000000001100110110100000; // input=-0.03564453125, output=1.60644841029
			11'd1061: out = 32'b00000000000000001100110111000000; // input=-0.03662109375, output=1.60742561094
			11'd1062: out = 32'b00000000000000001100110111100000; // input=-0.03759765625, output=1.60840284659
			11'd1063: out = 32'b00000000000000001100111000000000; // input=-0.03857421875, output=1.60938011817
			11'd1064: out = 32'b00000000000000001100111000100000; // input=-0.03955078125, output=1.61035742662
			11'd1065: out = 32'b00000000000000001100111001000000; // input=-0.04052734375, output=1.61133477288
			11'd1066: out = 32'b00000000000000001100111001100000; // input=-0.04150390625, output=1.61231215788
			11'd1067: out = 32'b00000000000000001100111010000000; // input=-0.04248046875, output=1.61328958257
			11'd1068: out = 32'b00000000000000001100111010100000; // input=-0.04345703125, output=1.61426704788
			11'd1069: out = 32'b00000000000000001100111011000000; // input=-0.04443359375, output=1.61524455475
			11'd1070: out = 32'b00000000000000001100111011100000; // input=-0.04541015625, output=1.61622210412
			11'd1071: out = 32'b00000000000000001100111100000000; // input=-0.04638671875, output=1.61719969694
			11'd1072: out = 32'b00000000000000001100111100100000; // input=-0.04736328125, output=1.61817733413
			11'd1073: out = 32'b00000000000000001100111101000000; // input=-0.04833984375, output=1.61915501665
			11'd1074: out = 32'b00000000000000001100111101100001; // input=-0.04931640625, output=1.62013274543
			11'd1075: out = 32'b00000000000000001100111110000001; // input=-0.05029296875, output=1.62111052141
			11'd1076: out = 32'b00000000000000001100111110100001; // input=-0.05126953125, output=1.62208834554
			11'd1077: out = 32'b00000000000000001100111111000001; // input=-0.05224609375, output=1.62306621875
			11'd1078: out = 32'b00000000000000001100111111100001; // input=-0.05322265625, output=1.624044142
			11'd1079: out = 32'b00000000000000001101000000000001; // input=-0.05419921875, output=1.62502211622
			11'd1080: out = 32'b00000000000000001101000000100001; // input=-0.05517578125, output=1.62600014235
			11'd1081: out = 32'b00000000000000001101000001000001; // input=-0.05615234375, output=1.62697822135
			11'd1082: out = 32'b00000000000000001101000001100001; // input=-0.05712890625, output=1.62795635416
			11'd1083: out = 32'b00000000000000001101000010000001; // input=-0.05810546875, output=1.62893454171
			11'd1084: out = 32'b00000000000000001101000010100001; // input=-0.05908203125, output=1.62991278496
			11'd1085: out = 32'b00000000000000001101000011000001; // input=-0.06005859375, output=1.63089108485
			11'd1086: out = 32'b00000000000000001101000011100001; // input=-0.06103515625, output=1.63186944233
			11'd1087: out = 32'b00000000000000001101000100000001; // input=-0.06201171875, output=1.63284785834
			11'd1088: out = 32'b00000000000000001101000100100001; // input=-0.06298828125, output=1.63382633383
			11'd1089: out = 32'b00000000000000001101000101000001; // input=-0.06396484375, output=1.63480486976
			11'd1090: out = 32'b00000000000000001101000101100001; // input=-0.06494140625, output=1.63578346706
			11'd1091: out = 32'b00000000000000001101000110000001; // input=-0.06591796875, output=1.63676212669
			11'd1092: out = 32'b00000000000000001101000110100001; // input=-0.06689453125, output=1.63774084959
			11'd1093: out = 32'b00000000000000001101000111000010; // input=-0.06787109375, output=1.63871963672
			11'd1094: out = 32'b00000000000000001101000111100010; // input=-0.06884765625, output=1.63969848903
			11'd1095: out = 32'b00000000000000001101001000000010; // input=-0.06982421875, output=1.64067740747
			11'd1096: out = 32'b00000000000000001101001000100010; // input=-0.07080078125, output=1.64165639298
			11'd1097: out = 32'b00000000000000001101001001000010; // input=-0.07177734375, output=1.64263544653
			11'd1098: out = 32'b00000000000000001101001001100010; // input=-0.07275390625, output=1.64361456906
			11'd1099: out = 32'b00000000000000001101001010000010; // input=-0.07373046875, output=1.64459376153
			11'd1100: out = 32'b00000000000000001101001010100010; // input=-0.07470703125, output=1.6455730249
			11'd1101: out = 32'b00000000000000001101001011000010; // input=-0.07568359375, output=1.64655236011
			11'd1102: out = 32'b00000000000000001101001011100010; // input=-0.07666015625, output=1.64753176812
			11'd1103: out = 32'b00000000000000001101001100000010; // input=-0.07763671875, output=1.64851124989
			11'd1104: out = 32'b00000000000000001101001100100011; // input=-0.07861328125, output=1.64949080637
			11'd1105: out = 32'b00000000000000001101001101000011; // input=-0.07958984375, output=1.65047043853
			11'd1106: out = 32'b00000000000000001101001101100011; // input=-0.08056640625, output=1.65145014731
			11'd1107: out = 32'b00000000000000001101001110000011; // input=-0.08154296875, output=1.65242993369
			11'd1108: out = 32'b00000000000000001101001110100011; // input=-0.08251953125, output=1.65340979861
			11'd1109: out = 32'b00000000000000001101001111000011; // input=-0.08349609375, output=1.65438974304
			11'd1110: out = 32'b00000000000000001101001111100011; // input=-0.08447265625, output=1.65536976794
			11'd1111: out = 32'b00000000000000001101010000000011; // input=-0.08544921875, output=1.65634987426
			11'd1112: out = 32'b00000000000000001101010000100011; // input=-0.08642578125, output=1.65733006298
			11'd1113: out = 32'b00000000000000001101010001000100; // input=-0.08740234375, output=1.65831033506
			11'd1114: out = 32'b00000000000000001101010001100100; // input=-0.08837890625, output=1.65929069145
			11'd1115: out = 32'b00000000000000001101010010000100; // input=-0.08935546875, output=1.66027113312
			11'd1116: out = 32'b00000000000000001101010010100100; // input=-0.09033203125, output=1.66125166104
			11'd1117: out = 32'b00000000000000001101010011000100; // input=-0.09130859375, output=1.66223227617
			11'd1118: out = 32'b00000000000000001101010011100100; // input=-0.09228515625, output=1.66321297948
			11'd1119: out = 32'b00000000000000001101010100000100; // input=-0.09326171875, output=1.66419377194
			11'd1120: out = 32'b00000000000000001101010100100100; // input=-0.09423828125, output=1.66517465451
			11'd1121: out = 32'b00000000000000001101010101000101; // input=-0.09521484375, output=1.66615562817
			11'd1122: out = 32'b00000000000000001101010101100101; // input=-0.09619140625, output=1.66713669388
			11'd1123: out = 32'b00000000000000001101010110000101; // input=-0.09716796875, output=1.66811785261
			11'd1124: out = 32'b00000000000000001101010110100101; // input=-0.09814453125, output=1.66909910534
			11'd1125: out = 32'b00000000000000001101010111000101; // input=-0.09912109375, output=1.67008045303
			11'd1126: out = 32'b00000000000000001101010111100101; // input=-0.10009765625, output=1.67106189666
			11'd1127: out = 32'b00000000000000001101011000000110; // input=-0.10107421875, output=1.67204343721
			11'd1128: out = 32'b00000000000000001101011000100110; // input=-0.10205078125, output=1.67302507565
			11'd1129: out = 32'b00000000000000001101011001000110; // input=-0.10302734375, output=1.67400681295
			11'd1130: out = 32'b00000000000000001101011001100110; // input=-0.10400390625, output=1.67498865008
			11'd1131: out = 32'b00000000000000001101011010000110; // input=-0.10498046875, output=1.67597058804
			11'd1132: out = 32'b00000000000000001101011010100110; // input=-0.10595703125, output=1.67695262779
			11'd1133: out = 32'b00000000000000001101011011000111; // input=-0.10693359375, output=1.67793477032
			11'd1134: out = 32'b00000000000000001101011011100111; // input=-0.10791015625, output=1.6789170166
			11'd1135: out = 32'b00000000000000001101011100000111; // input=-0.10888671875, output=1.67989936762
			11'd1136: out = 32'b00000000000000001101011100100111; // input=-0.10986328125, output=1.68088182435
			11'd1137: out = 32'b00000000000000001101011101000111; // input=-0.11083984375, output=1.68186438778
			11'd1138: out = 32'b00000000000000001101011101101000; // input=-0.11181640625, output=1.6828470589
			11'd1139: out = 32'b00000000000000001101011110001000; // input=-0.11279296875, output=1.68382983868
			11'd1140: out = 32'b00000000000000001101011110101000; // input=-0.11376953125, output=1.68481272812
			11'd1141: out = 32'b00000000000000001101011111001000; // input=-0.11474609375, output=1.6857957282
			11'd1142: out = 32'b00000000000000001101011111101000; // input=-0.11572265625, output=1.6867788399
			11'd1143: out = 32'b00000000000000001101100000001001; // input=-0.11669921875, output=1.68776206423
			11'd1144: out = 32'b00000000000000001101100000101001; // input=-0.11767578125, output=1.68874540215
			11'd1145: out = 32'b00000000000000001101100001001001; // input=-0.11865234375, output=1.68972885468
			11'd1146: out = 32'b00000000000000001101100001101001; // input=-0.11962890625, output=1.69071242279
			11'd1147: out = 32'b00000000000000001101100010001001; // input=-0.12060546875, output=1.69169610749
			11'd1148: out = 32'b00000000000000001101100010101010; // input=-0.12158203125, output=1.69267990976
			11'd1149: out = 32'b00000000000000001101100011001010; // input=-0.12255859375, output=1.69366383059
			11'd1150: out = 32'b00000000000000001101100011101010; // input=-0.12353515625, output=1.69464787099
			11'd1151: out = 32'b00000000000000001101100100001010; // input=-0.12451171875, output=1.69563203196
			11'd1152: out = 32'b00000000000000001101100100101011; // input=-0.12548828125, output=1.69661631448
			11'd1153: out = 32'b00000000000000001101100101001011; // input=-0.12646484375, output=1.69760071956
			11'd1154: out = 32'b00000000000000001101100101101011; // input=-0.12744140625, output=1.6985852482
			11'd1155: out = 32'b00000000000000001101100110001100; // input=-0.12841796875, output=1.69956990141
			11'd1156: out = 32'b00000000000000001101100110101100; // input=-0.12939453125, output=1.70055468017
			11'd1157: out = 32'b00000000000000001101100111001100; // input=-0.13037109375, output=1.7015395855
			11'd1158: out = 32'b00000000000000001101100111101100; // input=-0.13134765625, output=1.70252461839
			11'd1159: out = 32'b00000000000000001101101000001101; // input=-0.13232421875, output=1.70350977987
			11'd1160: out = 32'b00000000000000001101101000101101; // input=-0.13330078125, output=1.70449507093
			11'd1161: out = 32'b00000000000000001101101001001101; // input=-0.13427734375, output=1.70548049257
			11'd1162: out = 32'b00000000000000001101101001101101; // input=-0.13525390625, output=1.70646604582
			11'd1163: out = 32'b00000000000000001101101010001110; // input=-0.13623046875, output=1.70745173168
			11'd1164: out = 32'b00000000000000001101101010101110; // input=-0.13720703125, output=1.70843755116
			11'd1165: out = 32'b00000000000000001101101011001110; // input=-0.13818359375, output=1.70942350528
			11'd1166: out = 32'b00000000000000001101101011101111; // input=-0.13916015625, output=1.71040959504
			11'd1167: out = 32'b00000000000000001101101100001111; // input=-0.14013671875, output=1.71139582147
			11'd1168: out = 32'b00000000000000001101101100101111; // input=-0.14111328125, output=1.71238218558
			11'd1169: out = 32'b00000000000000001101101101010000; // input=-0.14208984375, output=1.71336868839
			11'd1170: out = 32'b00000000000000001101101101110000; // input=-0.14306640625, output=1.71435533091
			11'd1171: out = 32'b00000000000000001101101110010000; // input=-0.14404296875, output=1.71534211417
			11'd1172: out = 32'b00000000000000001101101110110001; // input=-0.14501953125, output=1.7163290392
			11'd1173: out = 32'b00000000000000001101101111010001; // input=-0.14599609375, output=1.717316107
			11'd1174: out = 32'b00000000000000001101101111110001; // input=-0.14697265625, output=1.71830331861
			11'd1175: out = 32'b00000000000000001101110000010010; // input=-0.14794921875, output=1.71929067505
			11'd1176: out = 32'b00000000000000001101110000110010; // input=-0.14892578125, output=1.72027817735
			11'd1177: out = 32'b00000000000000001101110001010010; // input=-0.14990234375, output=1.72126582653
			11'd1178: out = 32'b00000000000000001101110001110011; // input=-0.15087890625, output=1.72225362364
			11'd1179: out = 32'b00000000000000001101110010010011; // input=-0.15185546875, output=1.72324156968
			11'd1180: out = 32'b00000000000000001101110010110100; // input=-0.15283203125, output=1.72422966571
			11'd1181: out = 32'b00000000000000001101110011010100; // input=-0.15380859375, output=1.72521791275
			11'd1182: out = 32'b00000000000000001101110011110100; // input=-0.15478515625, output=1.72620631183
			11'd1183: out = 32'b00000000000000001101110100010101; // input=-0.15576171875, output=1.727194864
			11'd1184: out = 32'b00000000000000001101110100110101; // input=-0.15673828125, output=1.72818357029
			11'd1185: out = 32'b00000000000000001101110101010110; // input=-0.15771484375, output=1.72917243174
			11'd1186: out = 32'b00000000000000001101110101110110; // input=-0.15869140625, output=1.73016144939
			11'd1187: out = 32'b00000000000000001101110110010110; // input=-0.15966796875, output=1.73115062428
			11'd1188: out = 32'b00000000000000001101110110110111; // input=-0.16064453125, output=1.73213995746
			11'd1189: out = 32'b00000000000000001101110111010111; // input=-0.16162109375, output=1.73312944996
			11'd1190: out = 32'b00000000000000001101110111111000; // input=-0.16259765625, output=1.73411910285
			11'd1191: out = 32'b00000000000000001101111000011000; // input=-0.16357421875, output=1.73510891715
			11'd1192: out = 32'b00000000000000001101111000111000; // input=-0.16455078125, output=1.73609889394
			11'd1193: out = 32'b00000000000000001101111001011001; // input=-0.16552734375, output=1.73708903424
			11'd1194: out = 32'b00000000000000001101111001111001; // input=-0.16650390625, output=1.73807933913
			11'd1195: out = 32'b00000000000000001101111010011010; // input=-0.16748046875, output=1.73906980964
			11'd1196: out = 32'b00000000000000001101111010111010; // input=-0.16845703125, output=1.74006044684
			11'd1197: out = 32'b00000000000000001101111011011011; // input=-0.16943359375, output=1.74105125178
			11'd1198: out = 32'b00000000000000001101111011111011; // input=-0.17041015625, output=1.74204222552
			11'd1199: out = 32'b00000000000000001101111100011100; // input=-0.17138671875, output=1.74303336913
			11'd1200: out = 32'b00000000000000001101111100111100; // input=-0.17236328125, output=1.74402468365
			11'd1201: out = 32'b00000000000000001101111101011101; // input=-0.17333984375, output=1.74501617017
			11'd1202: out = 32'b00000000000000001101111101111101; // input=-0.17431640625, output=1.74600782973
			11'd1203: out = 32'b00000000000000001101111110011110; // input=-0.17529296875, output=1.74699966341
			11'd1204: out = 32'b00000000000000001101111110111110; // input=-0.17626953125, output=1.74799167227
			11'd1205: out = 32'b00000000000000001101111111011111; // input=-0.17724609375, output=1.74898385739
			11'd1206: out = 32'b00000000000000001101111111111111; // input=-0.17822265625, output=1.74997621983
			11'd1207: out = 32'b00000000000000001110000000100000; // input=-0.17919921875, output=1.75096876068
			11'd1208: out = 32'b00000000000000001110000001000000; // input=-0.18017578125, output=1.75196148099
			11'd1209: out = 32'b00000000000000001110000001100001; // input=-0.18115234375, output=1.75295438186
			11'd1210: out = 32'b00000000000000001110000010000001; // input=-0.18212890625, output=1.75394746435
			11'd1211: out = 32'b00000000000000001110000010100010; // input=-0.18310546875, output=1.75494072955
			11'd1212: out = 32'b00000000000000001110000011000010; // input=-0.18408203125, output=1.75593417853
			11'd1213: out = 32'b00000000000000001110000011100011; // input=-0.18505859375, output=1.75692781239
			11'd1214: out = 32'b00000000000000001110000100000100; // input=-0.18603515625, output=1.7579216322
			11'd1215: out = 32'b00000000000000001110000100100100; // input=-0.18701171875, output=1.75891563906
			11'd1216: out = 32'b00000000000000001110000101000101; // input=-0.18798828125, output=1.75990983405
			11'd1217: out = 32'b00000000000000001110000101100101; // input=-0.18896484375, output=1.76090421826
			11'd1218: out = 32'b00000000000000001110000110000110; // input=-0.18994140625, output=1.76189879278
			11'd1219: out = 32'b00000000000000001110000110100110; // input=-0.19091796875, output=1.76289355871
			11'd1220: out = 32'b00000000000000001110000111000111; // input=-0.19189453125, output=1.76388851714
			11'd1221: out = 32'b00000000000000001110000111101000; // input=-0.19287109375, output=1.76488366917
			11'd1222: out = 32'b00000000000000001110001000001000; // input=-0.19384765625, output=1.7658790159
			11'd1223: out = 32'b00000000000000001110001000101001; // input=-0.19482421875, output=1.76687455842
			11'd1224: out = 32'b00000000000000001110001001001010; // input=-0.19580078125, output=1.76787029786
			11'd1225: out = 32'b00000000000000001110001001101010; // input=-0.19677734375, output=1.76886623529
			11'd1226: out = 32'b00000000000000001110001010001011; // input=-0.19775390625, output=1.76986237185
			11'd1227: out = 32'b00000000000000001110001010101011; // input=-0.19873046875, output=1.77085870862
			11'd1228: out = 32'b00000000000000001110001011001100; // input=-0.19970703125, output=1.77185524673
			11'd1229: out = 32'b00000000000000001110001011101101; // input=-0.20068359375, output=1.77285198728
			11'd1230: out = 32'b00000000000000001110001100001101; // input=-0.20166015625, output=1.77384893139
			11'd1231: out = 32'b00000000000000001110001100101110; // input=-0.20263671875, output=1.77484608018
			11'd1232: out = 32'b00000000000000001110001101001111; // input=-0.20361328125, output=1.77584343476
			11'd1233: out = 32'b00000000000000001110001101110000; // input=-0.20458984375, output=1.77684099626
			11'd1234: out = 32'b00000000000000001110001110010000; // input=-0.20556640625, output=1.77783876579
			11'd1235: out = 32'b00000000000000001110001110110001; // input=-0.20654296875, output=1.77883674448
			11'd1236: out = 32'b00000000000000001110001111010010; // input=-0.20751953125, output=1.77983493346
			11'd1237: out = 32'b00000000000000001110001111110010; // input=-0.20849609375, output=1.78083333385
			11'd1238: out = 32'b00000000000000001110010000010011; // input=-0.20947265625, output=1.78183194679
			11'd1239: out = 32'b00000000000000001110010000110100; // input=-0.21044921875, output=1.78283077341
			11'd1240: out = 32'b00000000000000001110010001010101; // input=-0.21142578125, output=1.78382981483
			11'd1241: out = 32'b00000000000000001110010001110101; // input=-0.21240234375, output=1.78482907221
			11'd1242: out = 32'b00000000000000001110010010010110; // input=-0.21337890625, output=1.78582854667
			11'd1243: out = 32'b00000000000000001110010010110111; // input=-0.21435546875, output=1.78682823936
			11'd1244: out = 32'b00000000000000001110010011011000; // input=-0.21533203125, output=1.78782815142
			11'd1245: out = 32'b00000000000000001110010011111000; // input=-0.21630859375, output=1.788828284
			11'd1246: out = 32'b00000000000000001110010100011001; // input=-0.21728515625, output=1.78982863823
			11'd1247: out = 32'b00000000000000001110010100111010; // input=-0.21826171875, output=1.79082921528
			11'd1248: out = 32'b00000000000000001110010101011011; // input=-0.21923828125, output=1.79183001629
			11'd1249: out = 32'b00000000000000001110010101111011; // input=-0.22021484375, output=1.79283104241
			11'd1250: out = 32'b00000000000000001110010110011100; // input=-0.22119140625, output=1.79383229481
			11'd1251: out = 32'b00000000000000001110010110111101; // input=-0.22216796875, output=1.79483377464
			11'd1252: out = 32'b00000000000000001110010111011110; // input=-0.22314453125, output=1.79583548305
			11'd1253: out = 32'b00000000000000001110010111111111; // input=-0.22412109375, output=1.79683742122
			11'd1254: out = 32'b00000000000000001110011000100000; // input=-0.22509765625, output=1.79783959031
			11'd1255: out = 32'b00000000000000001110011001000000; // input=-0.22607421875, output=1.79884199148
			11'd1256: out = 32'b00000000000000001110011001100001; // input=-0.22705078125, output=1.7998446259
			11'd1257: out = 32'b00000000000000001110011010000010; // input=-0.22802734375, output=1.80084749474
			11'd1258: out = 32'b00000000000000001110011010100011; // input=-0.22900390625, output=1.80185059919
			11'd1259: out = 32'b00000000000000001110011011000100; // input=-0.22998046875, output=1.80285394041
			11'd1260: out = 32'b00000000000000001110011011100101; // input=-0.23095703125, output=1.80385751958
			11'd1261: out = 32'b00000000000000001110011100000110; // input=-0.23193359375, output=1.80486133789
			11'd1262: out = 32'b00000000000000001110011100100111; // input=-0.23291015625, output=1.80586539651
			11'd1263: out = 32'b00000000000000001110011101001000; // input=-0.23388671875, output=1.80686969664
			11'd1264: out = 32'b00000000000000001110011101101000; // input=-0.23486328125, output=1.80787423946
			11'd1265: out = 32'b00000000000000001110011110001001; // input=-0.23583984375, output=1.80887902616
			11'd1266: out = 32'b00000000000000001110011110101010; // input=-0.23681640625, output=1.80988405793
			11'd1267: out = 32'b00000000000000001110011111001011; // input=-0.23779296875, output=1.81088933598
			11'd1268: out = 32'b00000000000000001110011111101100; // input=-0.23876953125, output=1.81189486149
			11'd1269: out = 32'b00000000000000001110100000001101; // input=-0.23974609375, output=1.81290063567
			11'd1270: out = 32'b00000000000000001110100000101110; // input=-0.24072265625, output=1.81390665972
			11'd1271: out = 32'b00000000000000001110100001001111; // input=-0.24169921875, output=1.81491293484
			11'd1272: out = 32'b00000000000000001110100001110000; // input=-0.24267578125, output=1.81591946225
			11'd1273: out = 32'b00000000000000001110100010010001; // input=-0.24365234375, output=1.81692624315
			11'd1274: out = 32'b00000000000000001110100010110010; // input=-0.24462890625, output=1.81793327876
			11'd1275: out = 32'b00000000000000001110100011010011; // input=-0.24560546875, output=1.81894057029
			11'd1276: out = 32'b00000000000000001110100011110100; // input=-0.24658203125, output=1.81994811896
			11'd1277: out = 32'b00000000000000001110100100010101; // input=-0.24755859375, output=1.82095592599
			11'd1278: out = 32'b00000000000000001110100100110110; // input=-0.24853515625, output=1.82196399261
			11'd1279: out = 32'b00000000000000001110100101010111; // input=-0.24951171875, output=1.82297232004
			11'd1280: out = 32'b00000000000000001110100101111000; // input=-0.25048828125, output=1.8239809095
			11'd1281: out = 32'b00000000000000001110100110011001; // input=-0.25146484375, output=1.82498976223
			11'd1282: out = 32'b00000000000000001110100110111010; // input=-0.25244140625, output=1.82599887947
			11'd1283: out = 32'b00000000000000001110100111011011; // input=-0.25341796875, output=1.82700826245
			11'd1284: out = 32'b00000000000000001110100111111100; // input=-0.25439453125, output=1.82801791241
			11'd1285: out = 32'b00000000000000001110101000011110; // input=-0.25537109375, output=1.82902783059
			11'd1286: out = 32'b00000000000000001110101000111111; // input=-0.25634765625, output=1.83003801823
			11'd1287: out = 32'b00000000000000001110101001100000; // input=-0.25732421875, output=1.83104847659
			11'd1288: out = 32'b00000000000000001110101010000001; // input=-0.25830078125, output=1.83205920691
			11'd1289: out = 32'b00000000000000001110101010100010; // input=-0.25927734375, output=1.83307021045
			11'd1290: out = 32'b00000000000000001110101011000011; // input=-0.26025390625, output=1.83408148846
			11'd1291: out = 32'b00000000000000001110101011100100; // input=-0.26123046875, output=1.8350930422
			11'd1292: out = 32'b00000000000000001110101100000101; // input=-0.26220703125, output=1.83610487294
			11'd1293: out = 32'b00000000000000001110101100100111; // input=-0.26318359375, output=1.83711698194
			11'd1294: out = 32'b00000000000000001110101101001000; // input=-0.26416015625, output=1.83812937046
			11'd1295: out = 32'b00000000000000001110101101101001; // input=-0.26513671875, output=1.83914203977
			11'd1296: out = 32'b00000000000000001110101110001010; // input=-0.26611328125, output=1.84015499115
			11'd1297: out = 32'b00000000000000001110101110101011; // input=-0.26708984375, output=1.84116822588
			11'd1298: out = 32'b00000000000000001110101111001101; // input=-0.26806640625, output=1.84218174523
			11'd1299: out = 32'b00000000000000001110101111101110; // input=-0.26904296875, output=1.84319555049
			11'd1300: out = 32'b00000000000000001110110000001111; // input=-0.27001953125, output=1.84420964293
			11'd1301: out = 32'b00000000000000001110110000110000; // input=-0.27099609375, output=1.84522402386
			11'd1302: out = 32'b00000000000000001110110001010010; // input=-0.27197265625, output=1.84623869455
			11'd1303: out = 32'b00000000000000001110110001110011; // input=-0.27294921875, output=1.84725365631
			11'd1304: out = 32'b00000000000000001110110010010100; // input=-0.27392578125, output=1.84826891043
			11'd1305: out = 32'b00000000000000001110110010110101; // input=-0.27490234375, output=1.84928445821
			11'd1306: out = 32'b00000000000000001110110011010111; // input=-0.27587890625, output=1.85030030095
			11'd1307: out = 32'b00000000000000001110110011111000; // input=-0.27685546875, output=1.85131643996
			11'd1308: out = 32'b00000000000000001110110100011001; // input=-0.27783203125, output=1.85233287655
			11'd1309: out = 32'b00000000000000001110110100111011; // input=-0.27880859375, output=1.85334961204
			11'd1310: out = 32'b00000000000000001110110101011100; // input=-0.27978515625, output=1.85436664773
			11'd1311: out = 32'b00000000000000001110110101111101; // input=-0.28076171875, output=1.85538398495
			11'd1312: out = 32'b00000000000000001110110110011111; // input=-0.28173828125, output=1.85640162502
			11'd1313: out = 32'b00000000000000001110110111000000; // input=-0.28271484375, output=1.85741956927
			11'd1314: out = 32'b00000000000000001110110111100001; // input=-0.28369140625, output=1.85843781901
			11'd1315: out = 32'b00000000000000001110111000000011; // input=-0.28466796875, output=1.8594563756
			11'd1316: out = 32'b00000000000000001110111000100100; // input=-0.28564453125, output=1.86047524035
			11'd1317: out = 32'b00000000000000001110111001000101; // input=-0.28662109375, output=1.86149441461
			11'd1318: out = 32'b00000000000000001110111001100111; // input=-0.28759765625, output=1.86251389973
			11'd1319: out = 32'b00000000000000001110111010001000; // input=-0.28857421875, output=1.86353369704
			11'd1320: out = 32'b00000000000000001110111010101010; // input=-0.28955078125, output=1.86455380789
			11'd1321: out = 32'b00000000000000001110111011001011; // input=-0.29052734375, output=1.86557423364
			11'd1322: out = 32'b00000000000000001110111011101101; // input=-0.29150390625, output=1.86659497564
			11'd1323: out = 32'b00000000000000001110111100001110; // input=-0.29248046875, output=1.86761603526
			11'd1324: out = 32'b00000000000000001110111100110000; // input=-0.29345703125, output=1.86863741384
			11'd1325: out = 32'b00000000000000001110111101010001; // input=-0.29443359375, output=1.86965911277
			11'd1326: out = 32'b00000000000000001110111101110010; // input=-0.29541015625, output=1.8706811334
			11'd1327: out = 32'b00000000000000001110111110010100; // input=-0.29638671875, output=1.87170347712
			11'd1328: out = 32'b00000000000000001110111110110101; // input=-0.29736328125, output=1.87272614528
			11'd1329: out = 32'b00000000000000001110111111010111; // input=-0.29833984375, output=1.87374913929
			11'd1330: out = 32'b00000000000000001110111111111001; // input=-0.29931640625, output=1.87477246052
			11'd1331: out = 32'b00000000000000001111000000011010; // input=-0.30029296875, output=1.87579611035
			11'd1332: out = 32'b00000000000000001111000000111100; // input=-0.30126953125, output=1.87682009017
			11'd1333: out = 32'b00000000000000001111000001011101; // input=-0.30224609375, output=1.87784440139
			11'd1334: out = 32'b00000000000000001111000001111111; // input=-0.30322265625, output=1.8788690454
			11'd1335: out = 32'b00000000000000001111000010100000; // input=-0.30419921875, output=1.87989402359
			11'd1336: out = 32'b00000000000000001111000011000010; // input=-0.30517578125, output=1.88091933739
			11'd1337: out = 32'b00000000000000001111000011100100; // input=-0.30615234375, output=1.88194498818
			11'd1338: out = 32'b00000000000000001111000100000101; // input=-0.30712890625, output=1.88297097739
			11'd1339: out = 32'b00000000000000001111000100100111; // input=-0.30810546875, output=1.88399730643
			11'd1340: out = 32'b00000000000000001111000101001000; // input=-0.30908203125, output=1.88502397673
			11'd1341: out = 32'b00000000000000001111000101101010; // input=-0.31005859375, output=1.8860509897
			11'd1342: out = 32'b00000000000000001111000110001100; // input=-0.31103515625, output=1.88707834678
			11'd1343: out = 32'b00000000000000001111000110101101; // input=-0.31201171875, output=1.88810604939
			11'd1344: out = 32'b00000000000000001111000111001111; // input=-0.31298828125, output=1.88913409898
			11'd1345: out = 32'b00000000000000001111000111110001; // input=-0.31396484375, output=1.89016249697
			11'd1346: out = 32'b00000000000000001111001000010011; // input=-0.31494140625, output=1.89119124482
			11'd1347: out = 32'b00000000000000001111001000110100; // input=-0.31591796875, output=1.89222034396
			11'd1348: out = 32'b00000000000000001111001001010110; // input=-0.31689453125, output=1.89324979586
			11'd1349: out = 32'b00000000000000001111001001111000; // input=-0.31787109375, output=1.89427960197
			11'd1350: out = 32'b00000000000000001111001010011010; // input=-0.31884765625, output=1.89530976374
			11'd1351: out = 32'b00000000000000001111001010111011; // input=-0.31982421875, output=1.89634028265
			11'd1352: out = 32'b00000000000000001111001011011101; // input=-0.32080078125, output=1.89737116015
			11'd1353: out = 32'b00000000000000001111001011111111; // input=-0.32177734375, output=1.89840239771
			11'd1354: out = 32'b00000000000000001111001100100001; // input=-0.32275390625, output=1.89943399682
			11'd1355: out = 32'b00000000000000001111001101000010; // input=-0.32373046875, output=1.90046595895
			11'd1356: out = 32'b00000000000000001111001101100100; // input=-0.32470703125, output=1.90149828559
			11'd1357: out = 32'b00000000000000001111001110000110; // input=-0.32568359375, output=1.90253097822
			11'd1358: out = 32'b00000000000000001111001110101000; // input=-0.32666015625, output=1.90356403834
			11'd1359: out = 32'b00000000000000001111001111001010; // input=-0.32763671875, output=1.90459746744
			11'd1360: out = 32'b00000000000000001111001111101100; // input=-0.32861328125, output=1.90563126703
			11'd1361: out = 32'b00000000000000001111010000001110; // input=-0.32958984375, output=1.9066654386
			11'd1362: out = 32'b00000000000000001111010000110000; // input=-0.33056640625, output=1.90769998367
			11'd1363: out = 32'b00000000000000001111010001010001; // input=-0.33154296875, output=1.90873490375
			11'd1364: out = 32'b00000000000000001111010001110011; // input=-0.33251953125, output=1.90977020035
			11'd1365: out = 32'b00000000000000001111010010010101; // input=-0.33349609375, output=1.91080587501
			11'd1366: out = 32'b00000000000000001111010010110111; // input=-0.33447265625, output=1.91184192924
			11'd1367: out = 32'b00000000000000001111010011011001; // input=-0.33544921875, output=1.91287836459
			11'd1368: out = 32'b00000000000000001111010011111011; // input=-0.33642578125, output=1.91391518257
			11'd1369: out = 32'b00000000000000001111010100011101; // input=-0.33740234375, output=1.91495238474
			11'd1370: out = 32'b00000000000000001111010100111111; // input=-0.33837890625, output=1.91598997263
			11'd1371: out = 32'b00000000000000001111010101100001; // input=-0.33935546875, output=1.9170279478
			11'd1372: out = 32'b00000000000000001111010110000011; // input=-0.34033203125, output=1.91806631181
			11'd1373: out = 32'b00000000000000001111010110100101; // input=-0.34130859375, output=1.9191050662
			11'd1374: out = 32'b00000000000000001111010111000111; // input=-0.34228515625, output=1.92014421254
			11'd1375: out = 32'b00000000000000001111010111101001; // input=-0.34326171875, output=1.9211837524
			11'd1376: out = 32'b00000000000000001111011000001011; // input=-0.34423828125, output=1.92222368735
			11'd1377: out = 32'b00000000000000001111011000101110; // input=-0.34521484375, output=1.92326401896
			11'd1378: out = 32'b00000000000000001111011001010000; // input=-0.34619140625, output=1.92430474883
			11'd1379: out = 32'b00000000000000001111011001110010; // input=-0.34716796875, output=1.92534587853
			11'd1380: out = 32'b00000000000000001111011010010100; // input=-0.34814453125, output=1.92638740965
			11'd1381: out = 32'b00000000000000001111011010110110; // input=-0.34912109375, output=1.9274293438
			11'd1382: out = 32'b00000000000000001111011011011000; // input=-0.35009765625, output=1.92847168257
			11'd1383: out = 32'b00000000000000001111011011111010; // input=-0.35107421875, output=1.92951442757
			11'd1384: out = 32'b00000000000000001111011100011101; // input=-0.35205078125, output=1.93055758041
			11'd1385: out = 32'b00000000000000001111011100111111; // input=-0.35302734375, output=1.9316011427
			11'd1386: out = 32'b00000000000000001111011101100001; // input=-0.35400390625, output=1.93264511606
			11'd1387: out = 32'b00000000000000001111011110000011; // input=-0.35498046875, output=1.93368950212
			11'd1388: out = 32'b00000000000000001111011110100101; // input=-0.35595703125, output=1.93473430252
			11'd1389: out = 32'b00000000000000001111011111001000; // input=-0.35693359375, output=1.93577951888
			11'd1390: out = 32'b00000000000000001111011111101010; // input=-0.35791015625, output=1.93682515284
			11'd1391: out = 32'b00000000000000001111100000001100; // input=-0.35888671875, output=1.93787120606
			11'd1392: out = 32'b00000000000000001111100000101110; // input=-0.35986328125, output=1.93891768017
			11'd1393: out = 32'b00000000000000001111100001010001; // input=-0.36083984375, output=1.93996457685
			11'd1394: out = 32'b00000000000000001111100001110011; // input=-0.36181640625, output=1.94101189774
			11'd1395: out = 32'b00000000000000001111100010010101; // input=-0.36279296875, output=1.94205964452
			11'd1396: out = 32'b00000000000000001111100010111000; // input=-0.36376953125, output=1.94310781886
			11'd1397: out = 32'b00000000000000001111100011011010; // input=-0.36474609375, output=1.94415642243
			11'd1398: out = 32'b00000000000000001111100011111100; // input=-0.36572265625, output=1.94520545691
			11'd1399: out = 32'b00000000000000001111100100011111; // input=-0.36669921875, output=1.946254924
			11'd1400: out = 32'b00000000000000001111100101000001; // input=-0.36767578125, output=1.94730482538
			11'd1401: out = 32'b00000000000000001111100101100100; // input=-0.36865234375, output=1.94835516276
			11'd1402: out = 32'b00000000000000001111100110000110; // input=-0.36962890625, output=1.94940593784
			11'd1403: out = 32'b00000000000000001111100110101001; // input=-0.37060546875, output=1.95045715233
			11'd1404: out = 32'b00000000000000001111100111001011; // input=-0.37158203125, output=1.95150880793
			11'd1405: out = 32'b00000000000000001111100111101110; // input=-0.37255859375, output=1.95256090639
			11'd1406: out = 32'b00000000000000001111101000010000; // input=-0.37353515625, output=1.95361344941
			11'd1407: out = 32'b00000000000000001111101000110011; // input=-0.37451171875, output=1.95466643873
			11'd1408: out = 32'b00000000000000001111101001010101; // input=-0.37548828125, output=1.95571987608
			11'd1409: out = 32'b00000000000000001111101001111000; // input=-0.37646484375, output=1.95677376322
			11'd1410: out = 32'b00000000000000001111101010011010; // input=-0.37744140625, output=1.95782810189
			11'd1411: out = 32'b00000000000000001111101010111101; // input=-0.37841796875, output=1.95888289384
			11'd1412: out = 32'b00000000000000001111101011011111; // input=-0.37939453125, output=1.95993814083
			11'd1413: out = 32'b00000000000000001111101100000010; // input=-0.38037109375, output=1.96099384464
			11'd1414: out = 32'b00000000000000001111101100100100; // input=-0.38134765625, output=1.96205000703
			11'd1415: out = 32'b00000000000000001111101101000111; // input=-0.38232421875, output=1.96310662977
			11'd1416: out = 32'b00000000000000001111101101101010; // input=-0.38330078125, output=1.96416371466
			11'd1417: out = 32'b00000000000000001111101110001100; // input=-0.38427734375, output=1.96522126348
			11'd1418: out = 32'b00000000000000001111101110101111; // input=-0.38525390625, output=1.96627927804
			11'd1419: out = 32'b00000000000000001111101111010010; // input=-0.38623046875, output=1.96733776012
			11'd1420: out = 32'b00000000000000001111101111110100; // input=-0.38720703125, output=1.96839671154
			11'd1421: out = 32'b00000000000000001111110000010111; // input=-0.38818359375, output=1.96945613411
			11'd1422: out = 32'b00000000000000001111110000111010; // input=-0.38916015625, output=1.97051602965
			11'd1423: out = 32'b00000000000000001111110001011101; // input=-0.39013671875, output=1.9715764
			11'd1424: out = 32'b00000000000000001111110001111111; // input=-0.39111328125, output=1.97263724697
			11'd1425: out = 32'b00000000000000001111110010100010; // input=-0.39208984375, output=1.97369857241
			11'd1426: out = 32'b00000000000000001111110011000101; // input=-0.39306640625, output=1.97476037817
			11'd1427: out = 32'b00000000000000001111110011101000; // input=-0.39404296875, output=1.9758226661
			11'd1428: out = 32'b00000000000000001111110100001011; // input=-0.39501953125, output=1.97688543805
			11'd1429: out = 32'b00000000000000001111110100101101; // input=-0.39599609375, output=1.97794869588
			11'd1430: out = 32'b00000000000000001111110101010000; // input=-0.39697265625, output=1.97901244148
			11'd1431: out = 32'b00000000000000001111110101110011; // input=-0.39794921875, output=1.98007667672
			11'd1432: out = 32'b00000000000000001111110110010110; // input=-0.39892578125, output=1.98114140347
			11'd1433: out = 32'b00000000000000001111110110111001; // input=-0.39990234375, output=1.98220662364
			11'd1434: out = 32'b00000000000000001111110111011100; // input=-0.40087890625, output=1.98327233911
			11'd1435: out = 32'b00000000000000001111110111111111; // input=-0.40185546875, output=1.98433855179
			11'd1436: out = 32'b00000000000000001111111000100010; // input=-0.40283203125, output=1.9854052636
			11'd1437: out = 32'b00000000000000001111111001000101; // input=-0.40380859375, output=1.98647247644
			11'd1438: out = 32'b00000000000000001111111001101000; // input=-0.40478515625, output=1.98754019225
			11'd1439: out = 32'b00000000000000001111111010001011; // input=-0.40576171875, output=1.98860841295
			11'd1440: out = 32'b00000000000000001111111010101110; // input=-0.40673828125, output=1.98967714048
			11'd1441: out = 32'b00000000000000001111111011010001; // input=-0.40771484375, output=1.99074637679
			11'd1442: out = 32'b00000000000000001111111011110100; // input=-0.40869140625, output=1.99181612382
			11'd1443: out = 32'b00000000000000001111111100010111; // input=-0.40966796875, output=1.99288638354
			11'd1444: out = 32'b00000000000000001111111100111010; // input=-0.41064453125, output=1.99395715791
			11'd1445: out = 32'b00000000000000001111111101011101; // input=-0.41162109375, output=1.9950284489
			11'd1446: out = 32'b00000000000000001111111110000000; // input=-0.41259765625, output=1.9961002585
			11'd1447: out = 32'b00000000000000001111111110100011; // input=-0.41357421875, output=1.99717258869
			11'd1448: out = 32'b00000000000000001111111111000111; // input=-0.41455078125, output=1.99824544146
			11'd1449: out = 32'b00000000000000001111111111101010; // input=-0.41552734375, output=1.99931881882
			11'd1450: out = 32'b00000000000000010000000000001101; // input=-0.41650390625, output=2.00039272277
			11'd1451: out = 32'b00000000000000010000000000110000; // input=-0.41748046875, output=2.00146715533
			11'd1452: out = 32'b00000000000000010000000001010011; // input=-0.41845703125, output=2.00254211853
			11'd1453: out = 32'b00000000000000010000000001110111; // input=-0.41943359375, output=2.00361761439
			11'd1454: out = 32'b00000000000000010000000010011010; // input=-0.42041015625, output=2.00469364496
			11'd1455: out = 32'b00000000000000010000000010111101; // input=-0.42138671875, output=2.00577021228
			11'd1456: out = 32'b00000000000000010000000011100000; // input=-0.42236328125, output=2.0068473184
			11'd1457: out = 32'b00000000000000010000000100000100; // input=-0.42333984375, output=2.00792496538
			11'd1458: out = 32'b00000000000000010000000100100111; // input=-0.42431640625, output=2.0090031553
			11'd1459: out = 32'b00000000000000010000000101001010; // input=-0.42529296875, output=2.01008189023
			11'd1460: out = 32'b00000000000000010000000101101110; // input=-0.42626953125, output=2.01116117226
			11'd1461: out = 32'b00000000000000010000000110010001; // input=-0.42724609375, output=2.01224100347
			11'd1462: out = 32'b00000000000000010000000110110101; // input=-0.42822265625, output=2.01332138597
			11'd1463: out = 32'b00000000000000010000000111011000; // input=-0.42919921875, output=2.01440232187
			11'd1464: out = 32'b00000000000000010000000111111011; // input=-0.43017578125, output=2.01548381328
			11'd1465: out = 32'b00000000000000010000001000011111; // input=-0.43115234375, output=2.01656586232
			11'd1466: out = 32'b00000000000000010000001001000010; // input=-0.43212890625, output=2.01764847113
			11'd1467: out = 32'b00000000000000010000001001100110; // input=-0.43310546875, output=2.01873164186
			11'd1468: out = 32'b00000000000000010000001010001001; // input=-0.43408203125, output=2.01981537664
			11'd1469: out = 32'b00000000000000010000001010101101; // input=-0.43505859375, output=2.02089967763
			11'd1470: out = 32'b00000000000000010000001011010000; // input=-0.43603515625, output=2.02198454701
			11'd1471: out = 32'b00000000000000010000001011110100; // input=-0.43701171875, output=2.02306998694
			11'd1472: out = 32'b00000000000000010000001100011000; // input=-0.43798828125, output=2.0241559996
			11'd1473: out = 32'b00000000000000010000001100111011; // input=-0.43896484375, output=2.02524258719
			11'd1474: out = 32'b00000000000000010000001101011111; // input=-0.43994140625, output=2.02632975191
			11'd1475: out = 32'b00000000000000010000001110000010; // input=-0.44091796875, output=2.02741749596
			11'd1476: out = 32'b00000000000000010000001110100110; // input=-0.44189453125, output=2.02850582155
			11'd1477: out = 32'b00000000000000010000001111001010; // input=-0.44287109375, output=2.02959473092
			11'd1478: out = 32'b00000000000000010000001111101101; // input=-0.44384765625, output=2.0306842263
			11'd1479: out = 32'b00000000000000010000010000010001; // input=-0.44482421875, output=2.03177430993
			11'd1480: out = 32'b00000000000000010000010000110101; // input=-0.44580078125, output=2.03286498406
			11'd1481: out = 32'b00000000000000010000010001011001; // input=-0.44677734375, output=2.03395625095
			11'd1482: out = 32'b00000000000000010000010001111100; // input=-0.44775390625, output=2.03504811287
			11'd1483: out = 32'b00000000000000010000010010100000; // input=-0.44873046875, output=2.0361405721
			11'd1484: out = 32'b00000000000000010000010011000100; // input=-0.44970703125, output=2.03723363093
			11'd1485: out = 32'b00000000000000010000010011101000; // input=-0.45068359375, output=2.03832729165
			11'd1486: out = 32'b00000000000000010000010100001100; // input=-0.45166015625, output=2.03942155657
			11'd1487: out = 32'b00000000000000010000010100110000; // input=-0.45263671875, output=2.040516428
			11'd1488: out = 32'b00000000000000010000010101010100; // input=-0.45361328125, output=2.04161190827
			11'd1489: out = 32'b00000000000000010000010101110111; // input=-0.45458984375, output=2.0427079997
			11'd1490: out = 32'b00000000000000010000010110011011; // input=-0.45556640625, output=2.04380470466
			11'd1491: out = 32'b00000000000000010000010110111111; // input=-0.45654296875, output=2.04490202548
			11'd1492: out = 32'b00000000000000010000010111100011; // input=-0.45751953125, output=2.04599996453
			11'd1493: out = 32'b00000000000000010000011000000111; // input=-0.45849609375, output=2.04709852418
			11'd1494: out = 32'b00000000000000010000011000101011; // input=-0.45947265625, output=2.04819770681
			11'd1495: out = 32'b00000000000000010000011001001111; // input=-0.46044921875, output=2.04929751482
			11'd1496: out = 32'b00000000000000010000011001110011; // input=-0.46142578125, output=2.0503979506
			11'd1497: out = 32'b00000000000000010000011010011000; // input=-0.46240234375, output=2.05149901657
			11'd1498: out = 32'b00000000000000010000011010111100; // input=-0.46337890625, output=2.05260071515
			11'd1499: out = 32'b00000000000000010000011011100000; // input=-0.46435546875, output=2.05370304877
			11'd1500: out = 32'b00000000000000010000011100000100; // input=-0.46533203125, output=2.05480601986
			11'd1501: out = 32'b00000000000000010000011100101000; // input=-0.46630859375, output=2.05590963089
			11'd1502: out = 32'b00000000000000010000011101001100; // input=-0.46728515625, output=2.05701388431
			11'd1503: out = 32'b00000000000000010000011101110000; // input=-0.46826171875, output=2.05811878259
			11'd1504: out = 32'b00000000000000010000011110010101; // input=-0.46923828125, output=2.05922432822
			11'd1505: out = 32'b00000000000000010000011110111001; // input=-0.47021484375, output=2.0603305237
			11'd1506: out = 32'b00000000000000010000011111011101; // input=-0.47119140625, output=2.06143737151
			11'd1507: out = 32'b00000000000000010000100000000001; // input=-0.47216796875, output=2.06254487418
			11'd1508: out = 32'b00000000000000010000100000100110; // input=-0.47314453125, output=2.06365303424
			11'd1509: out = 32'b00000000000000010000100001001010; // input=-0.47412109375, output=2.06476185421
			11'd1510: out = 32'b00000000000000010000100001101110; // input=-0.47509765625, output=2.06587133664
			11'd1511: out = 32'b00000000000000010000100010010011; // input=-0.47607421875, output=2.06698148409
			11'd1512: out = 32'b00000000000000010000100010110111; // input=-0.47705078125, output=2.06809229913
			11'd1513: out = 32'b00000000000000010000100011011100; // input=-0.47802734375, output=2.06920378434
			11'd1514: out = 32'b00000000000000010000100100000000; // input=-0.47900390625, output=2.0703159423
			11'd1515: out = 32'b00000000000000010000100100100101; // input=-0.47998046875, output=2.07142877563
			11'd1516: out = 32'b00000000000000010000100101001001; // input=-0.48095703125, output=2.07254228692
			11'd1517: out = 32'b00000000000000010000100101101110; // input=-0.48193359375, output=2.07365647881
			11'd1518: out = 32'b00000000000000010000100110010010; // input=-0.48291015625, output=2.07477135392
			11'd1519: out = 32'b00000000000000010000100110110111; // input=-0.48388671875, output=2.07588691492
			11'd1520: out = 32'b00000000000000010000100111011011; // input=-0.48486328125, output=2.07700316444
			11'd1521: out = 32'b00000000000000010000101000000000; // input=-0.48583984375, output=2.07812010518
			11'd1522: out = 32'b00000000000000010000101000100100; // input=-0.48681640625, output=2.07923773979
			11'd1523: out = 32'b00000000000000010000101001001001; // input=-0.48779296875, output=2.08035607099
			11'd1524: out = 32'b00000000000000010000101001101110; // input=-0.48876953125, output=2.08147510147
			11'd1525: out = 32'b00000000000000010000101010010010; // input=-0.48974609375, output=2.08259483396
			11'd1526: out = 32'b00000000000000010000101010110111; // input=-0.49072265625, output=2.08371527118
			11'd1527: out = 32'b00000000000000010000101011011100; // input=-0.49169921875, output=2.08483641586
			11'd1528: out = 32'b00000000000000010000101100000001; // input=-0.49267578125, output=2.08595827078
			11'd1529: out = 32'b00000000000000010000101100100101; // input=-0.49365234375, output=2.08708083869
			11'd1530: out = 32'b00000000000000010000101101001010; // input=-0.49462890625, output=2.08820412237
			11'd1531: out = 32'b00000000000000010000101101101111; // input=-0.49560546875, output=2.08932812462
			11'd1532: out = 32'b00000000000000010000101110010100; // input=-0.49658203125, output=2.09045284823
			11'd1533: out = 32'b00000000000000010000101110111001; // input=-0.49755859375, output=2.09157829602
			11'd1534: out = 32'b00000000000000010000101111011110; // input=-0.49853515625, output=2.09270447082
			11'd1535: out = 32'b00000000000000010000110000000011; // input=-0.49951171875, output=2.09383137548
			11'd1536: out = 32'b00000000000000010000110000101000; // input=-0.50048828125, output=2.09495901284
			11'd1537: out = 32'b00000000000000010000110001001101; // input=-0.50146484375, output=2.09608738578
			11'd1538: out = 32'b00000000000000010000110001110010; // input=-0.50244140625, output=2.09721649718
			11'd1539: out = 32'b00000000000000010000110010010111; // input=-0.50341796875, output=2.09834634992
			11'd1540: out = 32'b00000000000000010000110010111100; // input=-0.50439453125, output=2.09947694693
			11'd1541: out = 32'b00000000000000010000110011100001; // input=-0.50537109375, output=2.10060829111
			11'd1542: out = 32'b00000000000000010000110100000110; // input=-0.50634765625, output=2.1017403854
			11'd1543: out = 32'b00000000000000010000110100101011; // input=-0.50732421875, output=2.10287323276
			11'd1544: out = 32'b00000000000000010000110101010000; // input=-0.50830078125, output=2.10400683614
			11'd1545: out = 32'b00000000000000010000110101110101; // input=-0.50927734375, output=2.10514119851
			11'd1546: out = 32'b00000000000000010000110110011010; // input=-0.51025390625, output=2.10627632287
			11'd1547: out = 32'b00000000000000010000110111000000; // input=-0.51123046875, output=2.10741221223
			11'd1548: out = 32'b00000000000000010000110111100101; // input=-0.51220703125, output=2.10854886959
			11'd1549: out = 32'b00000000000000010000111000001010; // input=-0.51318359375, output=2.10968629798
			11'd1550: out = 32'b00000000000000010000111000101111; // input=-0.51416015625, output=2.11082450046
			11'd1551: out = 32'b00000000000000010000111001010101; // input=-0.51513671875, output=2.11196348009
			11'd1552: out = 32'b00000000000000010000111001111010; // input=-0.51611328125, output=2.11310323994
			11'd1553: out = 32'b00000000000000010000111010100000; // input=-0.51708984375, output=2.11424378309
			11'd1554: out = 32'b00000000000000010000111011000101; // input=-0.51806640625, output=2.11538511266
			11'd1555: out = 32'b00000000000000010000111011101010; // input=-0.51904296875, output=2.11652723175
			11'd1556: out = 32'b00000000000000010000111100010000; // input=-0.52001953125, output=2.11767014351
			11'd1557: out = 32'b00000000000000010000111100110101; // input=-0.52099609375, output=2.11881385109
			11'd1558: out = 32'b00000000000000010000111101011011; // input=-0.52197265625, output=2.11995835764
			11'd1559: out = 32'b00000000000000010000111110000000; // input=-0.52294921875, output=2.12110366635
			11'd1560: out = 32'b00000000000000010000111110100110; // input=-0.52392578125, output=2.12224978041
			11'd1561: out = 32'b00000000000000010000111111001011; // input=-0.52490234375, output=2.12339670303
			11'd1562: out = 32'b00000000000000010000111111110001; // input=-0.52587890625, output=2.12454443744
			11'd1563: out = 32'b00000000000000010001000000010111; // input=-0.52685546875, output=2.12569298688
			11'd1564: out = 32'b00000000000000010001000000111100; // input=-0.52783203125, output=2.1268423546
			11'd1565: out = 32'b00000000000000010001000001100010; // input=-0.52880859375, output=2.12799254388
			11'd1566: out = 32'b00000000000000010001000010001000; // input=-0.52978515625, output=2.12914355801
			11'd1567: out = 32'b00000000000000010001000010101110; // input=-0.53076171875, output=2.13029540029
			11'd1568: out = 32'b00000000000000010001000011010011; // input=-0.53173828125, output=2.13144807404
			11'd1569: out = 32'b00000000000000010001000011111001; // input=-0.53271484375, output=2.13260158261
			11'd1570: out = 32'b00000000000000010001000100011111; // input=-0.53369140625, output=2.13375592934
			11'd1571: out = 32'b00000000000000010001000101000101; // input=-0.53466796875, output=2.13491111761
			11'd1572: out = 32'b00000000000000010001000101101011; // input=-0.53564453125, output=2.13606715081
			11'd1573: out = 32'b00000000000000010001000110010001; // input=-0.53662109375, output=2.13722403234
			11'd1574: out = 32'b00000000000000010001000110110110; // input=-0.53759765625, output=2.13838176562
			11'd1575: out = 32'b00000000000000010001000111011100; // input=-0.53857421875, output=2.1395403541
			11'd1576: out = 32'b00000000000000010001001000000010; // input=-0.53955078125, output=2.14069980123
			11'd1577: out = 32'b00000000000000010001001000101000; // input=-0.54052734375, output=2.14186011048
			11'd1578: out = 32'b00000000000000010001001001001111; // input=-0.54150390625, output=2.14302128534
			11'd1579: out = 32'b00000000000000010001001001110101; // input=-0.54248046875, output=2.14418332933
			11'd1580: out = 32'b00000000000000010001001010011011; // input=-0.54345703125, output=2.14534624597
			11'd1581: out = 32'b00000000000000010001001011000001; // input=-0.54443359375, output=2.14651003881
			11'd1582: out = 32'b00000000000000010001001011100111; // input=-0.54541015625, output=2.14767471141
			11'd1583: out = 32'b00000000000000010001001100001101; // input=-0.54638671875, output=2.14884026735
			11'd1584: out = 32'b00000000000000010001001100110011; // input=-0.54736328125, output=2.15000671023
			11'd1585: out = 32'b00000000000000010001001101011010; // input=-0.54833984375, output=2.15117404367
			11'd1586: out = 32'b00000000000000010001001110000000; // input=-0.54931640625, output=2.15234227131
			11'd1587: out = 32'b00000000000000010001001110100110; // input=-0.55029296875, output=2.1535113968
			11'd1588: out = 32'b00000000000000010001001111001101; // input=-0.55126953125, output=2.15468142383
			11'd1589: out = 32'b00000000000000010001001111110011; // input=-0.55224609375, output=2.15585235607
			11'd1590: out = 32'b00000000000000010001010000011001; // input=-0.55322265625, output=2.15702419726
			11'd1591: out = 32'b00000000000000010001010001000000; // input=-0.55419921875, output=2.15819695111
			11'd1592: out = 32'b00000000000000010001010001100110; // input=-0.55517578125, output=2.15937062138
			11'd1593: out = 32'b00000000000000010001010010001101; // input=-0.55615234375, output=2.16054521185
			11'd1594: out = 32'b00000000000000010001010010110011; // input=-0.55712890625, output=2.1617207263
			11'd1595: out = 32'b00000000000000010001010011011010; // input=-0.55810546875, output=2.16289716856
			11'd1596: out = 32'b00000000000000010001010100000000; // input=-0.55908203125, output=2.16407454244
			11'd1597: out = 32'b00000000000000010001010100100111; // input=-0.56005859375, output=2.16525285181
			11'd1598: out = 32'b00000000000000010001010101001110; // input=-0.56103515625, output=2.16643210053
			11'd1599: out = 32'b00000000000000010001010101110100; // input=-0.56201171875, output=2.16761229251
			11'd1600: out = 32'b00000000000000010001010110011011; // input=-0.56298828125, output=2.16879343165
			11'd1601: out = 32'b00000000000000010001010111000010; // input=-0.56396484375, output=2.1699755219
			11'd1602: out = 32'b00000000000000010001010111101001; // input=-0.56494140625, output=2.1711585672
			11'd1603: out = 32'b00000000000000010001011000001111; // input=-0.56591796875, output=2.17234257154
			11'd1604: out = 32'b00000000000000010001011000110110; // input=-0.56689453125, output=2.17352753892
			11'd1605: out = 32'b00000000000000010001011001011101; // input=-0.56787109375, output=2.17471347335
			11'd1606: out = 32'b00000000000000010001011010000100; // input=-0.56884765625, output=2.17590037889
			11'd1607: out = 32'b00000000000000010001011010101011; // input=-0.56982421875, output=2.1770882596
			11'd1608: out = 32'b00000000000000010001011011010010; // input=-0.57080078125, output=2.17827711957
			11'd1609: out = 32'b00000000000000010001011011111001; // input=-0.57177734375, output=2.1794669629
			11'd1610: out = 32'b00000000000000010001011100100000; // input=-0.57275390625, output=2.18065779373
			11'd1611: out = 32'b00000000000000010001011101000111; // input=-0.57373046875, output=2.18184961621
			11'd1612: out = 32'b00000000000000010001011101101110; // input=-0.57470703125, output=2.18304243453
			11'd1613: out = 32'b00000000000000010001011110010101; // input=-0.57568359375, output=2.18423625289
			11'd1614: out = 32'b00000000000000010001011110111100; // input=-0.57666015625, output=2.1854310755
			11'd1615: out = 32'b00000000000000010001011111100011; // input=-0.57763671875, output=2.18662690663
			11'd1616: out = 32'b00000000000000010001100000001011; // input=-0.57861328125, output=2.18782375054
			11'd1617: out = 32'b00000000000000010001100000110010; // input=-0.57958984375, output=2.18902161152
			11'd1618: out = 32'b00000000000000010001100001011001; // input=-0.58056640625, output=2.19022049391
			11'd1619: out = 32'b00000000000000010001100010000000; // input=-0.58154296875, output=2.19142040204
			11'd1620: out = 32'b00000000000000010001100010101000; // input=-0.58251953125, output=2.19262134028
			11'd1621: out = 32'b00000000000000010001100011001111; // input=-0.58349609375, output=2.19382331303
			11'd1622: out = 32'b00000000000000010001100011110111; // input=-0.58447265625, output=2.1950263247
			11'd1623: out = 32'b00000000000000010001100100011110; // input=-0.58544921875, output=2.19623037975
			11'd1624: out = 32'b00000000000000010001100101000110; // input=-0.58642578125, output=2.19743548264
			11'd1625: out = 32'b00000000000000010001100101101101; // input=-0.58740234375, output=2.19864163786
			11'd1626: out = 32'b00000000000000010001100110010101; // input=-0.58837890625, output=2.19984884994
			11'd1627: out = 32'b00000000000000010001100110111100; // input=-0.58935546875, output=2.20105712342
			11'd1628: out = 32'b00000000000000010001100111100100; // input=-0.59033203125, output=2.20226646288
			11'd1629: out = 32'b00000000000000010001101000001100; // input=-0.59130859375, output=2.20347687291
			11'd1630: out = 32'b00000000000000010001101000110011; // input=-0.59228515625, output=2.20468835815
			11'd1631: out = 32'b00000000000000010001101001011011; // input=-0.59326171875, output=2.20590092324
			11'd1632: out = 32'b00000000000000010001101010000011; // input=-0.59423828125, output=2.20711457287
			11'd1633: out = 32'b00000000000000010001101010101011; // input=-0.59521484375, output=2.20832931175
			11'd1634: out = 32'b00000000000000010001101011010010; // input=-0.59619140625, output=2.2095451446
			11'd1635: out = 32'b00000000000000010001101011111010; // input=-0.59716796875, output=2.21076207619
			11'd1636: out = 32'b00000000000000010001101100100010; // input=-0.59814453125, output=2.21198011132
			11'd1637: out = 32'b00000000000000010001101101001010; // input=-0.59912109375, output=2.21319925481
			11'd1638: out = 32'b00000000000000010001101101110010; // input=-0.60009765625, output=2.21441951149
			11'd1639: out = 32'b00000000000000010001101110011010; // input=-0.60107421875, output=2.21564088625
			11'd1640: out = 32'b00000000000000010001101111000010; // input=-0.60205078125, output=2.216863384
			11'd1641: out = 32'b00000000000000010001101111101010; // input=-0.60302734375, output=2.21808700967
			11'd1642: out = 32'b00000000000000010001110000010010; // input=-0.60400390625, output=2.21931176822
			11'd1643: out = 32'b00000000000000010001110000111011; // input=-0.60498046875, output=2.22053766465
			11'd1644: out = 32'b00000000000000010001110001100011; // input=-0.60595703125, output=2.22176470399
			11'd1645: out = 32'b00000000000000010001110010001011; // input=-0.60693359375, output=2.22299289128
			11'd1646: out = 32'b00000000000000010001110010110011; // input=-0.60791015625, output=2.22422223162
			11'd1647: out = 32'b00000000000000010001110011011100; // input=-0.60888671875, output=2.22545273013
			11'd1648: out = 32'b00000000000000010001110100000100; // input=-0.60986328125, output=2.22668439194
			11'd1649: out = 32'b00000000000000010001110100101100; // input=-0.61083984375, output=2.22791722224
			11'd1650: out = 32'b00000000000000010001110101010101; // input=-0.61181640625, output=2.22915122625
			11'd1651: out = 32'b00000000000000010001110101111101; // input=-0.61279296875, output=2.23038640919
			11'd1652: out = 32'b00000000000000010001110110100110; // input=-0.61376953125, output=2.23162277636
			11'd1653: out = 32'b00000000000000010001110111001110; // input=-0.61474609375, output=2.23286033305
			11'd1654: out = 32'b00000000000000010001110111110111; // input=-0.61572265625, output=2.23409908462
			11'd1655: out = 32'b00000000000000010001111000100000; // input=-0.61669921875, output=2.23533903642
			11'd1656: out = 32'b00000000000000010001111001001000; // input=-0.61767578125, output=2.23658019387
			11'd1657: out = 32'b00000000000000010001111001110001; // input=-0.61865234375, output=2.23782256242
			11'd1658: out = 32'b00000000000000010001111010011010; // input=-0.61962890625, output=2.23906614753
			11'd1659: out = 32'b00000000000000010001111011000011; // input=-0.62060546875, output=2.24031095471
			11'd1660: out = 32'b00000000000000010001111011101011; // input=-0.62158203125, output=2.24155698952
			11'd1661: out = 32'b00000000000000010001111100010100; // input=-0.62255859375, output=2.24280425753
			11'd1662: out = 32'b00000000000000010001111100111101; // input=-0.62353515625, output=2.24405276435
			11'd1663: out = 32'b00000000000000010001111101100110; // input=-0.62451171875, output=2.24530251564
			11'd1664: out = 32'b00000000000000010001111110001111; // input=-0.62548828125, output=2.24655351708
			11'd1665: out = 32'b00000000000000010001111110111000; // input=-0.62646484375, output=2.24780577439
			11'd1666: out = 32'b00000000000000010001111111100001; // input=-0.62744140625, output=2.24905929334
			11'd1667: out = 32'b00000000000000010010000000001010; // input=-0.62841796875, output=2.25031407972
			11'd1668: out = 32'b00000000000000010010000000110011; // input=-0.62939453125, output=2.25157013937
			11'd1669: out = 32'b00000000000000010010000001011101; // input=-0.63037109375, output=2.25282747815
			11'd1670: out = 32'b00000000000000010010000010000110; // input=-0.63134765625, output=2.25408610198
			11'd1671: out = 32'b00000000000000010010000010101111; // input=-0.63232421875, output=2.25534601681
			11'd1672: out = 32'b00000000000000010010000011011001; // input=-0.63330078125, output=2.25660722861
			11'd1673: out = 32'b00000000000000010010000100000010; // input=-0.63427734375, output=2.25786974343
			11'd1674: out = 32'b00000000000000010010000100101011; // input=-0.63525390625, output=2.25913356731
			11'd1675: out = 32'b00000000000000010010000101010101; // input=-0.63623046875, output=2.26039870638
			11'd1676: out = 32'b00000000000000010010000101111110; // input=-0.63720703125, output=2.26166516677
			11'd1677: out = 32'b00000000000000010010000110101000; // input=-0.63818359375, output=2.26293295467
			11'd1678: out = 32'b00000000000000010010000111010001; // input=-0.63916015625, output=2.26420207631
			11'd1679: out = 32'b00000000000000010010000111111011; // input=-0.64013671875, output=2.26547253796
			11'd1680: out = 32'b00000000000000010010001000100101; // input=-0.64111328125, output=2.26674434592
			11'd1681: out = 32'b00000000000000010010001001001110; // input=-0.64208984375, output=2.26801750655
			11'd1682: out = 32'b00000000000000010010001001111000; // input=-0.64306640625, output=2.26929202626
			11'd1683: out = 32'b00000000000000010010001010100010; // input=-0.64404296875, output=2.27056791146
			11'd1684: out = 32'b00000000000000010010001011001100; // input=-0.64501953125, output=2.27184516865
			11'd1685: out = 32'b00000000000000010010001011110110; // input=-0.64599609375, output=2.27312380436
			11'd1686: out = 32'b00000000000000010010001100100000; // input=-0.64697265625, output=2.27440382515
			11'd1687: out = 32'b00000000000000010010001101001010; // input=-0.64794921875, output=2.27568523764
			11'd1688: out = 32'b00000000000000010010001101110100; // input=-0.64892578125, output=2.27696804848
			11'd1689: out = 32'b00000000000000010010001110011110; // input=-0.64990234375, output=2.27825226439
			11'd1690: out = 32'b00000000000000010010001111001000; // input=-0.65087890625, output=2.27953789212
			11'd1691: out = 32'b00000000000000010010001111110010; // input=-0.65185546875, output=2.28082493846
			11'd1692: out = 32'b00000000000000010010010000011100; // input=-0.65283203125, output=2.28211341026
			11'd1693: out = 32'b00000000000000010010010001000111; // input=-0.65380859375, output=2.28340331442
			11'd1694: out = 32'b00000000000000010010010001110001; // input=-0.65478515625, output=2.28469465787
			11'd1695: out = 32'b00000000000000010010010010011011; // input=-0.65576171875, output=2.2859874476
			11'd1696: out = 32'b00000000000000010010010011000110; // input=-0.65673828125, output=2.28728169065
			11'd1697: out = 32'b00000000000000010010010011110000; // input=-0.65771484375, output=2.28857739412
			11'd1698: out = 32'b00000000000000010010010100011011; // input=-0.65869140625, output=2.28987456513
			11'd1699: out = 32'b00000000000000010010010101000101; // input=-0.65966796875, output=2.29117321088
			11'd1700: out = 32'b00000000000000010010010101110000; // input=-0.66064453125, output=2.2924733386
			11'd1701: out = 32'b00000000000000010010010110011010; // input=-0.66162109375, output=2.29377495559
			11'd1702: out = 32'b00000000000000010010010111000101; // input=-0.66259765625, output=2.29507806919
			11'd1703: out = 32'b00000000000000010010010111110000; // input=-0.66357421875, output=2.29638268678
			11'd1704: out = 32'b00000000000000010010011000011011; // input=-0.66455078125, output=2.29768881583
			11'd1705: out = 32'b00000000000000010010011001000110; // input=-0.66552734375, output=2.29899646382
			11'd1706: out = 32'b00000000000000010010011001110000; // input=-0.66650390625, output=2.30030563833
			11'd1707: out = 32'b00000000000000010010011010011011; // input=-0.66748046875, output=2.30161634695
			11'd1708: out = 32'b00000000000000010010011011000110; // input=-0.66845703125, output=2.30292859735
			11'd1709: out = 32'b00000000000000010010011011110001; // input=-0.66943359375, output=2.30424239726
			11'd1710: out = 32'b00000000000000010010011100011101; // input=-0.67041015625, output=2.30555775445
			11'd1711: out = 32'b00000000000000010010011101001000; // input=-0.67138671875, output=2.30687467675
			11'd1712: out = 32'b00000000000000010010011101110011; // input=-0.67236328125, output=2.30819317206
			11'd1713: out = 32'b00000000000000010010011110011110; // input=-0.67333984375, output=2.30951324833
			11'd1714: out = 32'b00000000000000010010011111001001; // input=-0.67431640625, output=2.31083491357
			11'd1715: out = 32'b00000000000000010010011111110101; // input=-0.67529296875, output=2.31215817585
			11'd1716: out = 32'b00000000000000010010100000100000; // input=-0.67626953125, output=2.3134830433
			11'd1717: out = 32'b00000000000000010010100001001100; // input=-0.67724609375, output=2.3148095241
			11'd1718: out = 32'b00000000000000010010100001110111; // input=-0.67822265625, output=2.3161376265
			11'd1719: out = 32'b00000000000000010010100010100011; // input=-0.67919921875, output=2.31746735883
			11'd1720: out = 32'b00000000000000010010100011001110; // input=-0.68017578125, output=2.31879872945
			11'd1721: out = 32'b00000000000000010010100011111010; // input=-0.68115234375, output=2.32013174681
			11'd1722: out = 32'b00000000000000010010100100100110; // input=-0.68212890625, output=2.3214664194
			11'd1723: out = 32'b00000000000000010010100101010010; // input=-0.68310546875, output=2.3228027558
			11'd1724: out = 32'b00000000000000010010100101111101; // input=-0.68408203125, output=2.32414076463
			11'd1725: out = 32'b00000000000000010010100110101001; // input=-0.68505859375, output=2.32548045461
			11'd1726: out = 32'b00000000000000010010100111010101; // input=-0.68603515625, output=2.32682183449
			11'd1727: out = 32'b00000000000000010010101000000001; // input=-0.68701171875, output=2.32816491311
			11'd1728: out = 32'b00000000000000010010101000101101; // input=-0.68798828125, output=2.32950969936
			11'd1729: out = 32'b00000000000000010010101001011001; // input=-0.68896484375, output=2.33085620223
			11'd1730: out = 32'b00000000000000010010101010000110; // input=-0.68994140625, output=2.33220443076
			11'd1731: out = 32'b00000000000000010010101010110010; // input=-0.69091796875, output=2.33355439404
			11'd1732: out = 32'b00000000000000010010101011011110; // input=-0.69189453125, output=2.33490610128
			11'd1733: out = 32'b00000000000000010010101100001011; // input=-0.69287109375, output=2.33625956172
			11'd1734: out = 32'b00000000000000010010101100110111; // input=-0.69384765625, output=2.33761478469
			11'd1735: out = 32'b00000000000000010010101101100011; // input=-0.69482421875, output=2.3389717796
			11'd1736: out = 32'b00000000000000010010101110010000; // input=-0.69580078125, output=2.34033055592
			11'd1737: out = 32'b00000000000000010010101110111101; // input=-0.69677734375, output=2.34169112321
			11'd1738: out = 32'b00000000000000010010101111101001; // input=-0.69775390625, output=2.34305349109
			11'd1739: out = 32'b00000000000000010010110000010110; // input=-0.69873046875, output=2.34441766927
			11'd1740: out = 32'b00000000000000010010110001000011; // input=-0.69970703125, output=2.34578366754
			11'd1741: out = 32'b00000000000000010010110001101111; // input=-0.70068359375, output=2.34715149575
			11'd1742: out = 32'b00000000000000010010110010011100; // input=-0.70166015625, output=2.34852116386
			11'd1743: out = 32'b00000000000000010010110011001001; // input=-0.70263671875, output=2.34989268189
			11'd1744: out = 32'b00000000000000010010110011110110; // input=-0.70361328125, output=2.35126605994
			11'd1745: out = 32'b00000000000000010010110100100011; // input=-0.70458984375, output=2.3526413082
			11'd1746: out = 32'b00000000000000010010110101010000; // input=-0.70556640625, output=2.35401843695
			11'd1747: out = 32'b00000000000000010010110101111110; // input=-0.70654296875, output=2.35539745654
			11'd1748: out = 32'b00000000000000010010110110101011; // input=-0.70751953125, output=2.35677837743
			11'd1749: out = 32'b00000000000000010010110111011000; // input=-0.70849609375, output=2.35816121012
			11'd1750: out = 32'b00000000000000010010111000000110; // input=-0.70947265625, output=2.35954596526
			11'd1751: out = 32'b00000000000000010010111000110011; // input=-0.71044921875, output=2.36093265353
			11'd1752: out = 32'b00000000000000010010111001100001; // input=-0.71142578125, output=2.36232128574
			11'd1753: out = 32'b00000000000000010010111010001110; // input=-0.71240234375, output=2.36371187278
			11'd1754: out = 32'b00000000000000010010111010111100; // input=-0.71337890625, output=2.36510442562
			11'd1755: out = 32'b00000000000000010010111011101001; // input=-0.71435546875, output=2.36649895534
			11'd1756: out = 32'b00000000000000010010111100010111; // input=-0.71533203125, output=2.36789547311
			11'd1757: out = 32'b00000000000000010010111101000101; // input=-0.71630859375, output=2.36929399018
			11'd1758: out = 32'b00000000000000010010111101110011; // input=-0.71728515625, output=2.37069451791
			11'd1759: out = 32'b00000000000000010010111110100001; // input=-0.71826171875, output=2.37209706777
			11'd1760: out = 32'b00000000000000010010111111001111; // input=-0.71923828125, output=2.3735016513
			11'd1761: out = 32'b00000000000000010010111111111101; // input=-0.72021484375, output=2.37490828016
			11'd1762: out = 32'b00000000000000010011000000101011; // input=-0.72119140625, output=2.37631696612
			11'd1763: out = 32'b00000000000000010011000001011001; // input=-0.72216796875, output=2.37772772102
			11'd1764: out = 32'b00000000000000010011000010001000; // input=-0.72314453125, output=2.37914055683
			11'd1765: out = 32'b00000000000000010011000010110110; // input=-0.72412109375, output=2.38055548562
			11'd1766: out = 32'b00000000000000010011000011100100; // input=-0.72509765625, output=2.38197251956
			11'd1767: out = 32'b00000000000000010011000100010011; // input=-0.72607421875, output=2.38339167094
			11'd1768: out = 32'b00000000000000010011000101000010; // input=-0.72705078125, output=2.38481295214
			11'd1769: out = 32'b00000000000000010011000101110000; // input=-0.72802734375, output=2.38623637568
			11'd1770: out = 32'b00000000000000010011000110011111; // input=-0.72900390625, output=2.38766195416
			11'd1771: out = 32'b00000000000000010011000111001110; // input=-0.72998046875, output=2.38908970031
			11'd1772: out = 32'b00000000000000010011000111111101; // input=-0.73095703125, output=2.39051962697
			11'd1773: out = 32'b00000000000000010011001000101011; // input=-0.73193359375, output=2.3919517471
			11'd1774: out = 32'b00000000000000010011001001011010; // input=-0.73291015625, output=2.39338607378
			11'd1775: out = 32'b00000000000000010011001010001010; // input=-0.73388671875, output=2.39482262021
			11'd1776: out = 32'b00000000000000010011001010111001; // input=-0.73486328125, output=2.39626139969
			11'd1777: out = 32'b00000000000000010011001011101000; // input=-0.73583984375, output=2.39770242567
			11'd1778: out = 32'b00000000000000010011001100010111; // input=-0.73681640625, output=2.39914571171
			11'd1779: out = 32'b00000000000000010011001101000111; // input=-0.73779296875, output=2.4005912715
			11'd1780: out = 32'b00000000000000010011001101110110; // input=-0.73876953125, output=2.40203911885
			11'd1781: out = 32'b00000000000000010011001110100110; // input=-0.73974609375, output=2.40348926771
			11'd1782: out = 32'b00000000000000010011001111010101; // input=-0.74072265625, output=2.40494173215
			11'd1783: out = 32'b00000000000000010011010000000101; // input=-0.74169921875, output=2.40639652638
			11'd1784: out = 32'b00000000000000010011010000110101; // input=-0.74267578125, output=2.40785366474
			11'd1785: out = 32'b00000000000000010011010001100100; // input=-0.74365234375, output=2.40931316171
			11'd1786: out = 32'b00000000000000010011010010010100; // input=-0.74462890625, output=2.4107750319
			11'd1787: out = 32'b00000000000000010011010011000100; // input=-0.74560546875, output=2.41223929006
			11'd1788: out = 32'b00000000000000010011010011110100; // input=-0.74658203125, output=2.4137059511
			11'd1789: out = 32'b00000000000000010011010100100100; // input=-0.74755859375, output=2.41517503004
			11'd1790: out = 32'b00000000000000010011010101010101; // input=-0.74853515625, output=2.41664654208
			11'd1791: out = 32'b00000000000000010011010110000101; // input=-0.74951171875, output=2.41812050255
			11'd1792: out = 32'b00000000000000010011010110110101; // input=-0.75048828125, output=2.41959692693
			11'd1793: out = 32'b00000000000000010011010111100110; // input=-0.75146484375, output=2.42107583084
			11'd1794: out = 32'b00000000000000010011011000010110; // input=-0.75244140625, output=2.42255723008
			11'd1795: out = 32'b00000000000000010011011001000111; // input=-0.75341796875, output=2.42404114058
			11'd1796: out = 32'b00000000000000010011011001111000; // input=-0.75439453125, output=2.42552757845
			11'd1797: out = 32'b00000000000000010011011010101000; // input=-0.75537109375, output=2.42701655995
			11'd1798: out = 32'b00000000000000010011011011011001; // input=-0.75634765625, output=2.42850810149
			11'd1799: out = 32'b00000000000000010011011100001010; // input=-0.75732421875, output=2.43000221966
			11'd1800: out = 32'b00000000000000010011011100111011; // input=-0.75830078125, output=2.43149893121
			11'd1801: out = 32'b00000000000000010011011101101100; // input=-0.75927734375, output=2.43299825307
			11'd1802: out = 32'b00000000000000010011011110011110; // input=-0.76025390625, output=2.43450020233
			11'd1803: out = 32'b00000000000000010011011111001111; // input=-0.76123046875, output=2.43600479626
			11'd1804: out = 32'b00000000000000010011100000000000; // input=-0.76220703125, output=2.4375120523
			11'd1805: out = 32'b00000000000000010011100000110010; // input=-0.76318359375, output=2.43902198807
			11'd1806: out = 32'b00000000000000010011100001100011; // input=-0.76416015625, output=2.44053462137
			11'd1807: out = 32'b00000000000000010011100010010101; // input=-0.76513671875, output=2.44204997021
			11'd1808: out = 32'b00000000000000010011100011000111; // input=-0.76611328125, output=2.44356805275
			11'd1809: out = 32'b00000000000000010011100011111001; // input=-0.76708984375, output=2.44508888736
			11'd1810: out = 32'b00000000000000010011100100101011; // input=-0.76806640625, output=2.44661249259
			11'd1811: out = 32'b00000000000000010011100101011101; // input=-0.76904296875, output=2.44813888721
			11'd1812: out = 32'b00000000000000010011100110001111; // input=-0.77001953125, output=2.44966809017
			11'd1813: out = 32'b00000000000000010011100111000001; // input=-0.77099609375, output=2.45120012061
			11'd1814: out = 32'b00000000000000010011100111110011; // input=-0.77197265625, output=2.4527349979
			11'd1815: out = 32'b00000000000000010011101000100110; // input=-0.77294921875, output=2.45427274161
			11'd1816: out = 32'b00000000000000010011101001011000; // input=-0.77392578125, output=2.4558133715
			11'd1817: out = 32'b00000000000000010011101010001011; // input=-0.77490234375, output=2.45735690757
			11'd1818: out = 32'b00000000000000010011101010111101; // input=-0.77587890625, output=2.45890337003
			11'd1819: out = 32'b00000000000000010011101011110000; // input=-0.77685546875, output=2.4604527793
			11'd1820: out = 32'b00000000000000010011101100100011; // input=-0.77783203125, output=2.46200515604
			11'd1821: out = 32'b00000000000000010011101101010110; // input=-0.77880859375, output=2.46356052112
			11'd1822: out = 32'b00000000000000010011101110001001; // input=-0.77978515625, output=2.46511889565
			11'd1823: out = 32'b00000000000000010011101110111100; // input=-0.78076171875, output=2.46668030098
			11'd1824: out = 32'b00000000000000010011101111101111; // input=-0.78173828125, output=2.46824475868
			11'd1825: out = 32'b00000000000000010011110000100011; // input=-0.78271484375, output=2.46981229058
			11'd1826: out = 32'b00000000000000010011110001010110; // input=-0.78369140625, output=2.47138291876
			11'd1827: out = 32'b00000000000000010011110010001010; // input=-0.78466796875, output=2.47295666552
			11'd1828: out = 32'b00000000000000010011110010111110; // input=-0.78564453125, output=2.47453355344
			11'd1829: out = 32'b00000000000000010011110011110001; // input=-0.78662109375, output=2.47611360534
			11'd1830: out = 32'b00000000000000010011110100100101; // input=-0.78759765625, output=2.47769684433
			11'd1831: out = 32'b00000000000000010011110101011001; // input=-0.78857421875, output=2.47928329375
			11'd1832: out = 32'b00000000000000010011110110001101; // input=-0.78955078125, output=2.48087297723
			11'd1833: out = 32'b00000000000000010011110111000001; // input=-0.79052734375, output=2.48246591868
			11'd1834: out = 32'b00000000000000010011110111110110; // input=-0.79150390625, output=2.48406214227
			11'd1835: out = 32'b00000000000000010011111000101010; // input=-0.79248046875, output=2.48566167247
			11'd1836: out = 32'b00000000000000010011111001011111; // input=-0.79345703125, output=2.48726453403
			11'd1837: out = 32'b00000000000000010011111010010011; // input=-0.79443359375, output=2.488870752
			11'd1838: out = 32'b00000000000000010011111011001000; // input=-0.79541015625, output=2.49048035171
			11'd1839: out = 32'b00000000000000010011111011111101; // input=-0.79638671875, output=2.49209335883
			11'd1840: out = 32'b00000000000000010011111100110010; // input=-0.79736328125, output=2.4937097993
			11'd1841: out = 32'b00000000000000010011111101100111; // input=-0.79833984375, output=2.49532969939
			11'd1842: out = 32'b00000000000000010011111110011100; // input=-0.79931640625, output=2.49695308569
			11'd1843: out = 32'b00000000000000010011111111010001; // input=-0.80029296875, output=2.49857998512
			11'd1844: out = 32'b00000000000000010100000000000111; // input=-0.80126953125, output=2.5002104249
			11'd1845: out = 32'b00000000000000010100000000111100; // input=-0.80224609375, output=2.50184443262
			11'd1846: out = 32'b00000000000000010100000001110010; // input=-0.80322265625, output=2.5034820362
			11'd1847: out = 32'b00000000000000010100000010101000; // input=-0.80419921875, output=2.50512326391
			11'd1848: out = 32'b00000000000000010100000011011110; // input=-0.80517578125, output=2.50676814435
			11'd1849: out = 32'b00000000000000010100000100010100; // input=-0.80615234375, output=2.50841670652
			11'd1850: out = 32'b00000000000000010100000101001010; // input=-0.80712890625, output=2.51006897974
			11'd1851: out = 32'b00000000000000010100000110000000; // input=-0.80810546875, output=2.51172499375
			11'd1852: out = 32'b00000000000000010100000110110111; // input=-0.80908203125, output=2.51338477864
			11'd1853: out = 32'b00000000000000010100000111101101; // input=-0.81005859375, output=2.51504836488
			11'd1854: out = 32'b00000000000000010100001000100100; // input=-0.81103515625, output=2.51671578336
			11'd1855: out = 32'b00000000000000010100001001011011; // input=-0.81201171875, output=2.51838706534
			11'd1856: out = 32'b00000000000000010100001010010001; // input=-0.81298828125, output=2.52006224252
			11'd1857: out = 32'b00000000000000010100001011001000; // input=-0.81396484375, output=2.52174134698
			11'd1858: out = 32'b00000000000000010100001100000000; // input=-0.81494140625, output=2.52342441124
			11'd1859: out = 32'b00000000000000010100001100110111; // input=-0.81591796875, output=2.52511146826
			11'd1860: out = 32'b00000000000000010100001101101110; // input=-0.81689453125, output=2.52680255142
			11'd1861: out = 32'b00000000000000010100001110100110; // input=-0.81787109375, output=2.52849769456
			11'd1862: out = 32'b00000000000000010100001111011101; // input=-0.81884765625, output=2.53019693197
			11'd1863: out = 32'b00000000000000010100010000010101; // input=-0.81982421875, output=2.53190029839
			11'd1864: out = 32'b00000000000000010100010001001101; // input=-0.82080078125, output=2.53360782906
			11'd1865: out = 32'b00000000000000010100010010000101; // input=-0.82177734375, output=2.53531955968
			11'd1866: out = 32'b00000000000000010100010010111110; // input=-0.82275390625, output=2.53703552645
			11'd1867: out = 32'b00000000000000010100010011110110; // input=-0.82373046875, output=2.53875576607
			11'd1868: out = 32'b00000000000000010100010100101110; // input=-0.82470703125, output=2.54048031574
			11'd1869: out = 32'b00000000000000010100010101100111; // input=-0.82568359375, output=2.54220921319
			11'd1870: out = 32'b00000000000000010100010110100000; // input=-0.82666015625, output=2.54394249668
			11'd1871: out = 32'b00000000000000010100010111011001; // input=-0.82763671875, output=2.54568020501
			11'd1872: out = 32'b00000000000000010100011000010010; // input=-0.82861328125, output=2.54742237753
			11'd1873: out = 32'b00000000000000010100011001001011; // input=-0.82958984375, output=2.54916905414
			11'd1874: out = 32'b00000000000000010100011010000101; // input=-0.83056640625, output=2.55092027535
			11'd1875: out = 32'b00000000000000010100011010111110; // input=-0.83154296875, output=2.55267608221
			11'd1876: out = 32'b00000000000000010100011011111000; // input=-0.83251953125, output=2.5544365164
			11'd1877: out = 32'b00000000000000010100011100110010; // input=-0.83349609375, output=2.55620162019
			11'd1878: out = 32'b00000000000000010100011101101100; // input=-0.83447265625, output=2.55797143649
			11'd1879: out = 32'b00000000000000010100011110100110; // input=-0.83544921875, output=2.55974600883
			11'd1880: out = 32'b00000000000000010100011111100000; // input=-0.83642578125, output=2.5615253814
			11'd1881: out = 32'b00000000000000010100100000011011; // input=-0.83740234375, output=2.56330959903
			11'd1882: out = 32'b00000000000000010100100001010101; // input=-0.83837890625, output=2.56509870727
			11'd1883: out = 32'b00000000000000010100100010010000; // input=-0.83935546875, output=2.5668927523
			11'd1884: out = 32'b00000000000000010100100011001011; // input=-0.84033203125, output=2.56869178106
			11'd1885: out = 32'b00000000000000010100100100000110; // input=-0.84130859375, output=2.57049584118
			11'd1886: out = 32'b00000000000000010100100101000001; // input=-0.84228515625, output=2.57230498103
			11'd1887: out = 32'b00000000000000010100100101111101; // input=-0.84326171875, output=2.57411924973
			11'd1888: out = 32'b00000000000000010100100110111000; // input=-0.84423828125, output=2.57593869719
			11'd1889: out = 32'b00000000000000010100100111110100; // input=-0.84521484375, output=2.57776337407
			11'd1890: out = 32'b00000000000000010100101000110000; // input=-0.84619140625, output=2.57959333186
			11'd1891: out = 32'b00000000000000010100101001101100; // input=-0.84716796875, output=2.58142862285
			11'd1892: out = 32'b00000000000000010100101010101001; // input=-0.84814453125, output=2.58326930019
			11'd1893: out = 32'b00000000000000010100101011100101; // input=-0.84912109375, output=2.58511541787
			11'd1894: out = 32'b00000000000000010100101100100010; // input=-0.85009765625, output=2.58696703077
			11'd1895: out = 32'b00000000000000010100101101011111; // input=-0.85107421875, output=2.58882419465
			11'd1896: out = 32'b00000000000000010100101110011100; // input=-0.85205078125, output=2.59068696621
			11'd1897: out = 32'b00000000000000010100101111011001; // input=-0.85302734375, output=2.59255540308
			11'd1898: out = 32'b00000000000000010100110000010110; // input=-0.85400390625, output=2.59442956385
			11'd1899: out = 32'b00000000000000010100110001010100; // input=-0.85498046875, output=2.59630950808
			11'd1900: out = 32'b00000000000000010100110010010010; // input=-0.85595703125, output=2.59819529636
			11'd1901: out = 32'b00000000000000010100110011010000; // input=-0.85693359375, output=2.60008699031
			11'd1902: out = 32'b00000000000000010100110100001110; // input=-0.85791015625, output=2.60198465258
			11'd1903: out = 32'b00000000000000010100110101001100; // input=-0.85888671875, output=2.60388834693
			11'd1904: out = 32'b00000000000000010100110110001011; // input=-0.85986328125, output=2.60579813822
			11'd1905: out = 32'b00000000000000010100110111001010; // input=-0.86083984375, output=2.60771409243
			11'd1906: out = 32'b00000000000000010100111000001001; // input=-0.86181640625, output=2.60963627672
			11'd1907: out = 32'b00000000000000010100111001001000; // input=-0.86279296875, output=2.61156475943
			11'd1908: out = 32'b00000000000000010100111010000111; // input=-0.86376953125, output=2.61349961013
			11'd1909: out = 32'b00000000000000010100111011000111; // input=-0.86474609375, output=2.61544089964
			11'd1910: out = 32'b00000000000000010100111100000111; // input=-0.86572265625, output=2.61738870006
			11'd1911: out = 32'b00000000000000010100111101000111; // input=-0.86669921875, output=2.61934308481
			11'd1912: out = 32'b00000000000000010100111110000111; // input=-0.86767578125, output=2.62130412866
			11'd1913: out = 32'b00000000000000010100111111000111; // input=-0.86865234375, output=2.62327190776
			11'd1914: out = 32'b00000000000000010101000000001000; // input=-0.86962890625, output=2.62524649969
			11'd1915: out = 32'b00000000000000010101000001001001; // input=-0.87060546875, output=2.62722798349
			11'd1916: out = 32'b00000000000000010101000010001010; // input=-0.87158203125, output=2.62921643969
			11'd1917: out = 32'b00000000000000010101000011001100; // input=-0.87255859375, output=2.63121195036
			11'd1918: out = 32'b00000000000000010101000100001101; // input=-0.87353515625, output=2.63321459915
			11'd1919: out = 32'b00000000000000010101000101001111; // input=-0.87451171875, output=2.63522447134
			11'd1920: out = 32'b00000000000000010101000110010001; // input=-0.87548828125, output=2.63724165386
			11'd1921: out = 32'b00000000000000010101000111010011; // input=-0.87646484375, output=2.63926623536
			11'd1922: out = 32'b00000000000000010101001000010110; // input=-0.87744140625, output=2.64129830626
			11'd1923: out = 32'b00000000000000010101001001011001; // input=-0.87841796875, output=2.64333795878
			11'd1924: out = 32'b00000000000000010101001010011100; // input=-0.87939453125, output=2.645385287
			11'd1925: out = 32'b00000000000000010101001011011111; // input=-0.88037109375, output=2.64744038691
			11'd1926: out = 32'b00000000000000010101001100100011; // input=-0.88134765625, output=2.64950335647
			11'd1927: out = 32'b00000000000000010101001101100111; // input=-0.88232421875, output=2.65157429567
			11'd1928: out = 32'b00000000000000010101001110101011; // input=-0.88330078125, output=2.65365330659
			11'd1929: out = 32'b00000000000000010101001111101111; // input=-0.88427734375, output=2.65574049343
			11'd1930: out = 32'b00000000000000010101010000110100; // input=-0.88525390625, output=2.65783596262
			11'd1931: out = 32'b00000000000000010101010001111001; // input=-0.88623046875, output=2.65993982287
			11'd1932: out = 32'b00000000000000010101010010111110; // input=-0.88720703125, output=2.66205218521
			11'd1933: out = 32'b00000000000000010101010100000100; // input=-0.88818359375, output=2.6641731631
			11'd1934: out = 32'b00000000000000010101010101001001; // input=-0.88916015625, output=2.66630287249
			11'd1935: out = 32'b00000000000000010101010110001111; // input=-0.89013671875, output=2.6684414319
			11'd1936: out = 32'b00000000000000010101010111010110; // input=-0.89111328125, output=2.67058896248
			11'd1937: out = 32'b00000000000000010101011000011101; // input=-0.89208984375, output=2.67274558811
			11'd1938: out = 32'b00000000000000010101011001100011; // input=-0.89306640625, output=2.67491143551
			11'd1939: out = 32'b00000000000000010101011010101011; // input=-0.89404296875, output=2.67708663428
			11'd1940: out = 32'b00000000000000010101011011110010; // input=-0.89501953125, output=2.67927131704
			11'd1941: out = 32'b00000000000000010101011100111010; // input=-0.89599609375, output=2.6814656195
			11'd1942: out = 32'b00000000000000010101011110000010; // input=-0.89697265625, output=2.68366968056
			11'd1943: out = 32'b00000000000000010101011111001011; // input=-0.89794921875, output=2.68588364245
			11'd1944: out = 32'b00000000000000010101100000010100; // input=-0.89892578125, output=2.6881076508
			11'd1945: out = 32'b00000000000000010101100001011101; // input=-0.89990234375, output=2.69034185478
			11'd1946: out = 32'b00000000000000010101100010100111; // input=-0.90087890625, output=2.69258640723
			11'd1947: out = 32'b00000000000000010101100011110001; // input=-0.90185546875, output=2.69484146476
			11'd1948: out = 32'b00000000000000010101100100111011; // input=-0.90283203125, output=2.69710718789
			11'd1949: out = 32'b00000000000000010101100110000101; // input=-0.90380859375, output=2.6993837412
			11'd1950: out = 32'b00000000000000010101100111010000; // input=-0.90478515625, output=2.70167129347
			11'd1951: out = 32'b00000000000000010101101000011100; // input=-0.90576171875, output=2.70397001782
			11'd1952: out = 32'b00000000000000010101101001100111; // input=-0.90673828125, output=2.70628009189
			11'd1953: out = 32'b00000000000000010101101010110011; // input=-0.90771484375, output=2.70860169798
			11'd1954: out = 32'b00000000000000010101101100000000; // input=-0.90869140625, output=2.71093502324
			11'd1955: out = 32'b00000000000000010101101101001101; // input=-0.90966796875, output=2.71328025987
			11'd1956: out = 32'b00000000000000010101101110011010; // input=-0.91064453125, output=2.71563760525
			11'd1957: out = 32'b00000000000000010101101111101000; // input=-0.91162109375, output=2.71800726222
			11'd1958: out = 32'b00000000000000010101110000110110; // input=-0.91259765625, output=2.72038943924
			11'd1959: out = 32'b00000000000000010101110010000100; // input=-0.91357421875, output=2.72278435059
			11'd1960: out = 32'b00000000000000010101110011010011; // input=-0.91455078125, output=2.72519221669
			11'd1961: out = 32'b00000000000000010101110100100010; // input=-0.91552734375, output=2.72761326425
			11'd1962: out = 32'b00000000000000010101110101110010; // input=-0.91650390625, output=2.73004772657
			11'd1963: out = 32'b00000000000000010101110111000010; // input=-0.91748046875, output=2.73249584383
			11'd1964: out = 32'b00000000000000010101111000010011; // input=-0.91845703125, output=2.73495786332
			11'd1965: out = 32'b00000000000000010101111001100100; // input=-0.91943359375, output=2.73743403981
			11'd1966: out = 32'b00000000000000010101111010110110; // input=-0.92041015625, output=2.73992463579
			11'd1967: out = 32'b00000000000000010101111100001000; // input=-0.92138671875, output=2.74242992187
			11'd1968: out = 32'b00000000000000010101111101011011; // input=-0.92236328125, output=2.74495017711
			11'd1969: out = 32'b00000000000000010101111110101110; // input=-0.92333984375, output=2.74748568938
			11'd1970: out = 32'b00000000000000010110000000000001; // input=-0.92431640625, output=2.75003675577
			11'd1971: out = 32'b00000000000000010110000001010101; // input=-0.92529296875, output=2.752603683
			11'd1972: out = 32'b00000000000000010110000010101010; // input=-0.92626953125, output=2.75518678789
			11'd1973: out = 32'b00000000000000010110000011111111; // input=-0.92724609375, output=2.75778639778
			11'd1974: out = 32'b00000000000000010110000101010101; // input=-0.92822265625, output=2.76040285107
			11'd1975: out = 32'b00000000000000010110000110101011; // input=-0.92919921875, output=2.76303649773
			11'd1976: out = 32'b00000000000000010110001000000010; // input=-0.93017578125, output=2.76568769986
			11'd1977: out = 32'b00000000000000010110001001011010; // input=-0.93115234375, output=2.76835683229
			11'd1978: out = 32'b00000000000000010110001010110010; // input=-0.93212890625, output=2.77104428323
			11'd1979: out = 32'b00000000000000010110001100001010; // input=-0.93310546875, output=2.77375045491
			11'd1980: out = 32'b00000000000000010110001101100100; // input=-0.93408203125, output=2.77647576435
			11'd1981: out = 32'b00000000000000010110001110111110; // input=-0.93505859375, output=2.77922064407
			11'd1982: out = 32'b00000000000000010110010000011000; // input=-0.93603515625, output=2.78198554298
			11'd1983: out = 32'b00000000000000010110010001110011; // input=-0.93701171875, output=2.7847709272
			11'd1984: out = 32'b00000000000000010110010011001111; // input=-0.93798828125, output=2.78757728101
			11'd1985: out = 32'b00000000000000010110010100101100; // input=-0.93896484375, output=2.79040510791
			11'd1986: out = 32'b00000000000000010110010110001001; // input=-0.93994140625, output=2.79325493161
			11'd1987: out = 32'b00000000000000010110010111100111; // input=-0.94091796875, output=2.79612729726
			11'd1988: out = 32'b00000000000000010110011001000110; // input=-0.94189453125, output=2.79902277268
			11'd1989: out = 32'b00000000000000010110011010100110; // input=-0.94287109375, output=2.80194194967
			11'd1990: out = 32'b00000000000000010110011100000110; // input=-0.94384765625, output=2.8048854455
			11'd1991: out = 32'b00000000000000010110011101101000; // input=-0.94482421875, output=2.80785390442
			11'd1992: out = 32'b00000000000000010110011111001010; // input=-0.94580078125, output=2.81084799938
			11'd1993: out = 32'b00000000000000010110100000101101; // input=-0.94677734375, output=2.81386843382
			11'd1994: out = 32'b00000000000000010110100010010001; // input=-0.94775390625, output=2.81691594366
			11'd1995: out = 32'b00000000000000010110100011110101; // input=-0.94873046875, output=2.81999129943
			11'd1996: out = 32'b00000000000000010110100101011011; // input=-0.94970703125, output=2.8230953086
			11'd1997: out = 32'b00000000000000010110100111000010; // input=-0.95068359375, output=2.82622881808
			11'd1998: out = 32'b00000000000000010110101000101010; // input=-0.95166015625, output=2.82939271698
			11'd1999: out = 32'b00000000000000010110101010010010; // input=-0.95263671875, output=2.83258793963
			11'd2000: out = 32'b00000000000000010110101011111100; // input=-0.95361328125, output=2.83581546885
			11'd2001: out = 32'b00000000000000010110101101100111; // input=-0.95458984375, output=2.83907633955
			11'd2002: out = 32'b00000000000000010110101111010011; // input=-0.95556640625, output=2.84237164265
			11'd2003: out = 32'b00000000000000010110110001000000; // input=-0.95654296875, output=2.84570252945
			11'd2004: out = 32'b00000000000000010110110010101110; // input=-0.95751953125, output=2.84907021641
			11'd2005: out = 32'b00000000000000010110110100011110; // input=-0.95849609375, output=2.85247599038
			11'd2006: out = 32'b00000000000000010110110110001111; // input=-0.95947265625, output=2.85592121451
			11'd2007: out = 32'b00000000000000010110111000000001; // input=-0.96044921875, output=2.85940733468
			11'd2008: out = 32'b00000000000000010110111001110101; // input=-0.96142578125, output=2.86293588669
			11'd2009: out = 32'b00000000000000010110111011101010; // input=-0.96240234375, output=2.86650850434
			11'd2010: out = 32'b00000000000000010110111101100000; // input=-0.96337890625, output=2.87012692836
			11'd2011: out = 32'b00000000000000010110111111011000; // input=-0.96435546875, output=2.87379301647
			11'd2012: out = 32'b00000000000000010111000001010010; // input=-0.96533203125, output=2.87750875471
			11'd2013: out = 32'b00000000000000010111000011001110; // input=-0.96630859375, output=2.88127627019
			11'd2014: out = 32'b00000000000000010111000101001011; // input=-0.96728515625, output=2.88509784549
			11'd2015: out = 32'b00000000000000010111000111001010; // input=-0.96826171875, output=2.88897593506
			11'd2016: out = 32'b00000000000000010111001001001011; // input=-0.96923828125, output=2.89291318391
			11'd2017: out = 32'b00000000000000010111001011001110; // input=-0.97021484375, output=2.89691244895
			11'd2018: out = 32'b00000000000000010111001101010011; // input=-0.97119140625, output=2.90097682353
			11'd2019: out = 32'b00000000000000010111001111011011; // input=-0.97216796875, output=2.90510966579
			11'd2020: out = 32'b00000000000000010111010001100100; // input=-0.97314453125, output=2.90931463147
			11'd2021: out = 32'b00000000000000010111010011110001; // input=-0.97412109375, output=2.91359571221
			11'd2022: out = 32'b00000000000000010111010110000000; // input=-0.97509765625, output=2.91795728034
			11'd2023: out = 32'b00000000000000010111011000010001; // input=-0.97607421875, output=2.92240414177
			11'd2024: out = 32'b00000000000000010111011010100110; // input=-0.97705078125, output=2.92694159862
			11'd2025: out = 32'b00000000000000010111011100111110; // input=-0.97802734375, output=2.93157552401
			11'd2026: out = 32'b00000000000000010111011111011001; // input=-0.97900390625, output=2.93631245203
			11'd2027: out = 32'b00000000000000010111100001111000; // input=-0.97998046875, output=2.94115968675
			11'd2028: out = 32'b00000000000000010111100100011011; // input=-0.98095703125, output=2.94612543553
			11'd2029: out = 32'b00000000000000010111100111000010; // input=-0.98193359375, output=2.95121897351
			11'd2030: out = 32'b00000000000000010111101001101101; // input=-0.98291015625, output=2.95645084881
			11'd2031: out = 32'b00000000000000010111101100011101; // input=-0.98388671875, output=2.9618331413
			11'd2032: out = 32'b00000000000000010111101111010011; // input=-0.98486328125, output=2.96737979326
			11'd2033: out = 32'b00000000000000010111110010001111; // input=-0.98583984375, output=2.97310703786
			11'd2034: out = 32'b00000000000000010111110101010001; // input=-0.98681640625, output=2.97903396338
			11'd2035: out = 32'b00000000000000010111111000011010; // input=-0.98779296875, output=2.98518326972
			11'd2036: out = 32'b00000000000000010111111011101100; // input=-0.98876953125, output=2.99158230393
			11'd2037: out = 32'b00000000000000010111111111000111; // input=-0.98974609375, output=2.99826451197
			11'd2038: out = 32'b00000000000000011000000010101101; // input=-0.99072265625, output=3.00527153127
			11'd2039: out = 32'b00000000000000011000000110011111; // input=-0.99169921875, output=3.01265630832
			11'd2040: out = 32'b00000000000000011000001010011111; // input=-0.99267578125, output=3.02048793072
			11'd2041: out = 32'b00000000000000011000001110110010; // input=-0.99365234375, output=3.0288594899
			11'd2042: out = 32'b00000000000000011000010011011010; // input=-0.99462890625, output=3.03790168237
			11'd2043: out = 32'b00000000000000011000011000011111; // input=-0.99560546875, output=3.04780828732
			11'd2044: out = 32'b00000000000000011000011110001010; // input=-0.99658203125, output=3.05888935726
			11'd2045: out = 32'b00000000000000011000100100101110; // input=-0.99755859375, output=3.07170130494
			11'd2046: out = 32'b00000000000000011000101100110010; // input=-0.99853515625, output=3.08745945643
			11'd2047: out = 32'b00000000000000011000111000100000; // input=-0.99951171875, output=3.11034138188
		endcase
	end
	converter U0 (a, index);

endmodule

module asin_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000000000000000010000; // input=0.00048828125, output=0.000488281269403
			11'd1: out = 32'b00000000000000000000000000110000; // input=0.00146484375, output=0.00146484427387
			11'd2: out = 32'b00000000000000000000000001010000; // input=0.00244140625, output=0.00244140867533
			11'd3: out = 32'b00000000000000000000000001110000; // input=0.00341796875, output=0.00341797540511
			11'd4: out = 32'b00000000000000000000000010010000; // input=0.00439453125, output=0.00439454539458
			11'd5: out = 32'b00000000000000000000000010110000; // input=0.00537109375, output=0.00537111957513
			11'd6: out = 32'b00000000000000000000000011010000; // input=0.00634765625, output=0.00634769887818
			11'd7: out = 32'b00000000000000000000000011110000; // input=0.00732421875, output=0.0073242842352
			11'd8: out = 32'b00000000000000000000000100010000; // input=0.00830078125, output=0.0083008765777
			11'd9: out = 32'b00000000000000000000000100110000; // input=0.00927734375, output=0.00927747683727
			11'd10: out = 32'b00000000000000000000000101010000; // input=0.01025390625, output=0.0102540859456
			11'd11: out = 32'b00000000000000000000000101110000; // input=0.01123046875, output=0.0112307048343
			11'd12: out = 32'b00000000000000000000000110010000; // input=0.01220703125, output=0.0122073344352
			11'd13: out = 32'b00000000000000000000000110110000; // input=0.01318359375, output=0.0131839756803
			11'd14: out = 32'b00000000000000000000000111010000; // input=0.01416015625, output=0.0141606295016
			11'd15: out = 32'b00000000000000000000000111110000; // input=0.01513671875, output=0.0151372968311
			11'd16: out = 32'b00000000000000000000001000010000; // input=0.01611328125, output=0.016113978601
			11'd17: out = 32'b00000000000000000000001000110000; // input=0.01708984375, output=0.0170906757438
			11'd18: out = 32'b00000000000000000000001001010000; // input=0.01806640625, output=0.0180673891919
			11'd19: out = 32'b00000000000000000000001001110000; // input=0.01904296875, output=0.0190441198779
			11'd20: out = 32'b00000000000000000000001010010000; // input=0.02001953125, output=0.0200208687346
			11'd21: out = 32'b00000000000000000000001010110000; // input=0.02099609375, output=0.0209976366949
			11'd22: out = 32'b00000000000000000000001011010000; // input=0.02197265625, output=0.0219744246919
			11'd23: out = 32'b00000000000000000000001011110000; // input=0.02294921875, output=0.0229512336589
			11'd24: out = 32'b00000000000000000000001100010000; // input=0.02392578125, output=0.0239280645293
			11'd25: out = 32'b00000000000000000000001100110000; // input=0.02490234375, output=0.0249049182366
			11'd26: out = 32'b00000000000000000000001101010000; // input=0.02587890625, output=0.0258817957149
			11'd27: out = 32'b00000000000000000000001101110000; // input=0.02685546875, output=0.026858697898
			11'd28: out = 32'b00000000000000000000001110010000; // input=0.02783203125, output=0.0278356257202
			11'd29: out = 32'b00000000000000000000001110110000; // input=0.02880859375, output=0.028812580116
			11'd30: out = 32'b00000000000000000000001111010000; // input=0.02978515625, output=0.0297895620201
			11'd31: out = 32'b00000000000000000000001111110000; // input=0.03076171875, output=0.0307665723674
			11'd32: out = 32'b00000000000000000000010000010000; // input=0.03173828125, output=0.0317436120931
			11'd33: out = 32'b00000000000000000000010000110000; // input=0.03271484375, output=0.0327206821325
			11'd34: out = 32'b00000000000000000000010001010000; // input=0.03369140625, output=0.0336977834215
			11'd35: out = 32'b00000000000000000000010001110000; // input=0.03466796875, output=0.0346749168959
			11'd36: out = 32'b00000000000000000000010010010000; // input=0.03564453125, output=0.0356520834919
			11'd37: out = 32'b00000000000000000000010010110000; // input=0.03662109375, output=0.0366292841462
			11'd38: out = 32'b00000000000000000000010011010000; // input=0.03759765625, output=0.0376065197954
			11'd39: out = 32'b00000000000000000000010011110000; // input=0.03857421875, output=0.0385837913767
			11'd40: out = 32'b00000000000000000000010100010000; // input=0.03955078125, output=0.0395610998276
			11'd41: out = 32'b00000000000000000000010100110000; // input=0.04052734375, output=0.0405384460857
			11'd42: out = 32'b00000000000000000000010101010000; // input=0.04150390625, output=0.0415158310892
			11'd43: out = 32'b00000000000000000000010101110000; // input=0.04248046875, output=0.0424932557764
			11'd44: out = 32'b00000000000000000000010110010000; // input=0.04345703125, output=0.0434707210861
			11'd45: out = 32'b00000000000000000000010110110000; // input=0.04443359375, output=0.0444482279573
			11'd46: out = 32'b00000000000000000000010111010001; // input=0.04541015625, output=0.0454257773296
			11'd47: out = 32'b00000000000000000000010111110001; // input=0.04638671875, output=0.0464033701426
			11'd48: out = 32'b00000000000000000000011000010001; // input=0.04736328125, output=0.0473810073367
			11'd49: out = 32'b00000000000000000000011000110001; // input=0.04833984375, output=0.0483586898524
			11'd50: out = 32'b00000000000000000000011001010001; // input=0.04931640625, output=0.0493364186307
			11'd51: out = 32'b00000000000000000000011001110001; // input=0.05029296875, output=0.0503141946129
			11'd52: out = 32'b00000000000000000000011010010001; // input=0.05126953125, output=0.0512920187407
			11'd53: out = 32'b00000000000000000000011010110001; // input=0.05224609375, output=0.0522698919565
			11'd54: out = 32'b00000000000000000000011011010001; // input=0.05322265625, output=0.0532478152028
			11'd55: out = 32'b00000000000000000000011011110001; // input=0.05419921875, output=0.0542257894226
			11'd56: out = 32'b00000000000000000000011100010001; // input=0.05517578125, output=0.0552038155595
			11'd57: out = 32'b00000000000000000000011100110001; // input=0.05615234375, output=0.0561818945573
			11'd58: out = 32'b00000000000000000000011101010001; // input=0.05712890625, output=0.0571600273605
			11'd59: out = 32'b00000000000000000000011101110001; // input=0.05810546875, output=0.0581382149139
			11'd60: out = 32'b00000000000000000000011110010001; // input=0.05908203125, output=0.0591164581629
			11'd61: out = 32'b00000000000000000000011110110001; // input=0.06005859375, output=0.0600947580532
			11'd62: out = 32'b00000000000000000000011111010001; // input=0.06103515625, output=0.0610731155313
			11'd63: out = 32'b00000000000000000000011111110001; // input=0.06201171875, output=0.0620515315438
			11'd64: out = 32'b00000000000000000000100000010001; // input=0.06298828125, output=0.0630300070381
			11'd65: out = 32'b00000000000000000000100000110001; // input=0.06396484375, output=0.064008542962
			11'd66: out = 32'b00000000000000000000100001010001; // input=0.06494140625, output=0.064987140264
			11'd67: out = 32'b00000000000000000000100001110010; // input=0.06591796875, output=0.0659657998927
			11'd68: out = 32'b00000000000000000000100010010010; // input=0.06689453125, output=0.0669445227978
			11'd69: out = 32'b00000000000000000000100010110010; // input=0.06787109375, output=0.0679233099292
			11'd70: out = 32'b00000000000000000000100011010010; // input=0.06884765625, output=0.0689021622373
			11'd71: out = 32'b00000000000000000000100011110010; // input=0.06982421875, output=0.0698810806733
			11'd72: out = 32'b00000000000000000000100100010010; // input=0.07080078125, output=0.070860066189
			11'd73: out = 32'b00000000000000000000100100110010; // input=0.07177734375, output=0.0718391197364
			11'd74: out = 32'b00000000000000000000100101010010; // input=0.07275390625, output=0.0728182422686
			11'd75: out = 32'b00000000000000000000100101110010; // input=0.07373046875, output=0.0737974347388
			11'd76: out = 32'b00000000000000000000100110010010; // input=0.07470703125, output=0.0747766981013
			11'd77: out = 32'b00000000000000000000100110110010; // input=0.07568359375, output=0.0757560333106
			11'd78: out = 32'b00000000000000000000100111010010; // input=0.07666015625, output=0.0767354413221
			11'd79: out = 32'b00000000000000000000100111110011; // input=0.07763671875, output=0.0777149230917
			11'd80: out = 32'b00000000000000000000101000010011; // input=0.07861328125, output=0.0786944795761
			11'd81: out = 32'b00000000000000000000101000110011; // input=0.07958984375, output=0.0796741117323
			11'd82: out = 32'b00000000000000000000101001010011; // input=0.08056640625, output=0.0806538205183
			11'd83: out = 32'b00000000000000000000101001110011; // input=0.08154296875, output=0.0816336068927
			11'd84: out = 32'b00000000000000000000101010010011; // input=0.08251953125, output=0.0826134718148
			11'd85: out = 32'b00000000000000000000101010110011; // input=0.08349609375, output=0.0835934162443
			11'd86: out = 32'b00000000000000000000101011010011; // input=0.08447265625, output=0.084573441142
			11'd87: out = 32'b00000000000000000000101011110011; // input=0.08544921875, output=0.0855535474692
			11'd88: out = 32'b00000000000000000000101100010100; // input=0.08642578125, output=0.086533736188
			11'd89: out = 32'b00000000000000000000101100110100; // input=0.08740234375, output=0.087514008261
			11'd90: out = 32'b00000000000000000000101101010100; // input=0.08837890625, output=0.0884943646517
			11'd91: out = 32'b00000000000000000000101101110100; // input=0.08935546875, output=0.0894748063244
			11'd92: out = 32'b00000000000000000000101110010100; // input=0.09033203125, output=0.0904553342441
			11'd93: out = 32'b00000000000000000000101110110100; // input=0.09130859375, output=0.0914359493765
			11'd94: out = 32'b00000000000000000000101111010100; // input=0.09228515625, output=0.0924166526881
			11'd95: out = 32'b00000000000000000000101111110100; // input=0.09326171875, output=0.0933974451461
			11'd96: out = 32'b00000000000000000000110000010101; // input=0.09423828125, output=0.0943783277186
			11'd97: out = 32'b00000000000000000000110000110101; // input=0.09521484375, output=0.0953593013745
			11'd98: out = 32'b00000000000000000000110001010101; // input=0.09619140625, output=0.0963403670833
			11'd99: out = 32'b00000000000000000000110001110101; // input=0.09716796875, output=0.0973215258156
			11'd100: out = 32'b00000000000000000000110010010101; // input=0.09814453125, output=0.0983027785426
			11'd101: out = 32'b00000000000000000000110010110101; // input=0.09912109375, output=0.0992841262364
			11'd102: out = 32'b00000000000000000000110011010110; // input=0.10009765625, output=0.10026556987
			11'd103: out = 32'b00000000000000000000110011110110; // input=0.10107421875, output=0.101247110417
			11'd104: out = 32'b00000000000000000000110100010110; // input=0.10205078125, output=0.102228748852
			11'd105: out = 32'b00000000000000000000110100110110; // input=0.10302734375, output=0.103210486151
			11'd106: out = 32'b00000000000000000000110101010110; // input=0.10400390625, output=0.10419232329
			11'd107: out = 32'b00000000000000000000110101110110; // input=0.10498046875, output=0.105174261246
			11'd108: out = 32'b00000000000000000000110110010111; // input=0.10595703125, output=0.106156300998
			11'd109: out = 32'b00000000000000000000110110110111; // input=0.10693359375, output=0.107138443524
			11'd110: out = 32'b00000000000000000000110111010111; // input=0.10791015625, output=0.108120689804
			11'd111: out = 32'b00000000000000000000110111110111; // input=0.10888671875, output=0.10910304082
			11'd112: out = 32'b00000000000000000000111000010111; // input=0.10986328125, output=0.110085497553
			11'd113: out = 32'b00000000000000000000111000110111; // input=0.11083984375, output=0.111068060986
			11'd114: out = 32'b00000000000000000000111001011000; // input=0.11181640625, output=0.112050732102
			11'd115: out = 32'b00000000000000000000111001111000; // input=0.11279296875, output=0.113033511886
			11'd116: out = 32'b00000000000000000000111010011000; // input=0.11376953125, output=0.114016401324
			11'd117: out = 32'b00000000000000000000111010111000; // input=0.11474609375, output=0.114999401402
			11'd118: out = 32'b00000000000000000000111011011001; // input=0.11572265625, output=0.115982513109
			11'd119: out = 32'b00000000000000000000111011111001; // input=0.11669921875, output=0.116965737431
			11'd120: out = 32'b00000000000000000000111100011001; // input=0.11767578125, output=0.11794907536
			11'd121: out = 32'b00000000000000000000111100111001; // input=0.11865234375, output=0.118932527885
			11'd122: out = 32'b00000000000000000000111101011001; // input=0.11962890625, output=0.119916095998
			11'd123: out = 32'b00000000000000000000111101111010; // input=0.12060546875, output=0.120899780692
			11'd124: out = 32'b00000000000000000000111110011010; // input=0.12158203125, output=0.12188358296
			11'd125: out = 32'b00000000000000000000111110111010; // input=0.12255859375, output=0.122867503798
			11'd126: out = 32'b00000000000000000000111111011010; // input=0.12353515625, output=0.1238515442
			11'd127: out = 32'b00000000000000000000111111111011; // input=0.12451171875, output=0.124835705164
			11'd128: out = 32'b00000000000000000001000000011011; // input=0.12548828125, output=0.125819987687
			11'd129: out = 32'b00000000000000000001000000111011; // input=0.12646484375, output=0.126804392769
			11'd130: out = 32'b00000000000000000001000001011011; // input=0.12744140625, output=0.12778892141
			11'd131: out = 32'b00000000000000000001000001111100; // input=0.12841796875, output=0.12877357461
			11'd132: out = 32'b00000000000000000001000010011100; // input=0.12939453125, output=0.129758353373
			11'd133: out = 32'b00000000000000000001000010111100; // input=0.13037109375, output=0.130743258701
			11'd134: out = 32'b00000000000000000001000011011100; // input=0.13134765625, output=0.1317282916
			11'd135: out = 32'b00000000000000000001000011111101; // input=0.13232421875, output=0.132713453074
			11'd136: out = 32'b00000000000000000001000100011101; // input=0.13330078125, output=0.133698744131
			11'd137: out = 32'b00000000000000000001000100111101; // input=0.13427734375, output=0.134684165779
			11'd138: out = 32'b00000000000000000001000101011110; // input=0.13525390625, output=0.135669719027
			11'd139: out = 32'b00000000000000000001000101111110; // input=0.13623046875, output=0.136655404886
			11'd140: out = 32'b00000000000000000001000110011110; // input=0.13720703125, output=0.137641224367
			11'd141: out = 32'b00000000000000000001000110111111; // input=0.13818359375, output=0.138627178482
			11'd142: out = 32'b00000000000000000001000111011111; // input=0.13916015625, output=0.139613268246
			11'd143: out = 32'b00000000000000000001000111111111; // input=0.14013671875, output=0.140599494675
			11'd144: out = 32'b00000000000000000001001000011111; // input=0.14111328125, output=0.141585858784
			11'd145: out = 32'b00000000000000000001001001000000; // input=0.14208984375, output=0.142572361592
			11'd146: out = 32'b00000000000000000001001001100000; // input=0.14306640625, output=0.143559004117
			11'd147: out = 32'b00000000000000000001001010000000; // input=0.14404296875, output=0.144545787379
			11'd148: out = 32'b00000000000000000001001010100001; // input=0.14501953125, output=0.145532712401
			11'd149: out = 32'b00000000000000000001001011000001; // input=0.14599609375, output=0.146519780204
			11'd150: out = 32'b00000000000000000001001011100010; // input=0.14697265625, output=0.147506991814
			11'd151: out = 32'b00000000000000000001001100000010; // input=0.14794921875, output=0.148494348255
			11'd152: out = 32'b00000000000000000001001100100010; // input=0.14892578125, output=0.149481850554
			11'd153: out = 32'b00000000000000000001001101000011; // input=0.14990234375, output=0.15046949974
			11'd154: out = 32'b00000000000000000001001101100011; // input=0.15087890625, output=0.151457296841
			11'd155: out = 32'b00000000000000000001001110000011; // input=0.15185546875, output=0.152445242889
			11'd156: out = 32'b00000000000000000001001110100100; // input=0.15283203125, output=0.153433338915
			11'd157: out = 32'b00000000000000000001001111000100; // input=0.15380859375, output=0.154421585953
			11'd158: out = 32'b00000000000000000001001111100100; // input=0.15478515625, output=0.155409985038
			11'd159: out = 32'b00000000000000000001010000000101; // input=0.15576171875, output=0.156398537206
			11'd160: out = 32'b00000000000000000001010000100101; // input=0.15673828125, output=0.157387243495
			11'd161: out = 32'b00000000000000000001010001000110; // input=0.15771484375, output=0.158376104944
			11'd162: out = 32'b00000000000000000001010001100110; // input=0.15869140625, output=0.159365122593
			11'd163: out = 32'b00000000000000000001010010000110; // input=0.15966796875, output=0.160354297484
			11'd164: out = 32'b00000000000000000001010010100111; // input=0.16064453125, output=0.161343630661
			11'd165: out = 32'b00000000000000000001010011000111; // input=0.16162109375, output=0.162333123168
			11'd166: out = 32'b00000000000000000001010011101000; // input=0.16259765625, output=0.163322776052
			11'd167: out = 32'b00000000000000000001010100001000; // input=0.16357421875, output=0.16431259036
			11'd168: out = 32'b00000000000000000001010100101001; // input=0.16455078125, output=0.165302567142
			11'd169: out = 32'b00000000000000000001010101001001; // input=0.16552734375, output=0.166292707448
			11'd170: out = 32'b00000000000000000001010101101010; // input=0.16650390625, output=0.167283012331
			11'd171: out = 32'b00000000000000000001010110001010; // input=0.16748046875, output=0.168273482845
			11'd172: out = 32'b00000000000000000001010110101010; // input=0.16845703125, output=0.169264120044
			11'd173: out = 32'b00000000000000000001010111001011; // input=0.16943359375, output=0.170254924986
			11'd174: out = 32'b00000000000000000001010111101011; // input=0.17041015625, output=0.171245898729
			11'd175: out = 32'b00000000000000000001011000001100; // input=0.17138671875, output=0.172237042333
			11'd176: out = 32'b00000000000000000001011000101100; // input=0.17236328125, output=0.173228356859
			11'd177: out = 32'b00000000000000000001011001001101; // input=0.17333984375, output=0.174219843372
			11'd178: out = 32'b00000000000000000001011001101101; // input=0.17431640625, output=0.175211502934
			11'd179: out = 32'b00000000000000000001011010001110; // input=0.17529296875, output=0.176203336613
			11'd180: out = 32'b00000000000000000001011010101110; // input=0.17626953125, output=0.177195345477
			11'd181: out = 32'b00000000000000000001011011001111; // input=0.17724609375, output=0.178187530595
			11'd182: out = 32'b00000000000000000001011011101111; // input=0.17822265625, output=0.179179893039
			11'd183: out = 32'b00000000000000000001011100010000; // input=0.17919921875, output=0.180172433881
			11'd184: out = 32'b00000000000000000001011100110000; // input=0.18017578125, output=0.181165154197
			11'd185: out = 32'b00000000000000000001011101010001; // input=0.18115234375, output=0.182158055061
			11'd186: out = 32'b00000000000000000001011101110001; // input=0.18212890625, output=0.183151137553
			11'd187: out = 32'b00000000000000000001011110010010; // input=0.18310546875, output=0.184144402751
			11'd188: out = 32'b00000000000000000001011110110011; // input=0.18408203125, output=0.185137851738
			11'd189: out = 32'b00000000000000000001011111010011; // input=0.18505859375, output=0.186131485596
			11'd190: out = 32'b00000000000000000001011111110100; // input=0.18603515625, output=0.187125305409
			11'd191: out = 32'b00000000000000000001100000010100; // input=0.18701171875, output=0.188119312266
			11'd192: out = 32'b00000000000000000001100000110101; // input=0.18798828125, output=0.189113507254
			11'd193: out = 32'b00000000000000000001100001010101; // input=0.18896484375, output=0.190107891462
			11'd194: out = 32'b00000000000000000001100001110110; // input=0.18994140625, output=0.191102465984
			11'd195: out = 32'b00000000000000000001100010010111; // input=0.19091796875, output=0.192097231912
			11'd196: out = 32'b00000000000000000001100010110111; // input=0.19189453125, output=0.193092190343
			11'd197: out = 32'b00000000000000000001100011011000; // input=0.19287109375, output=0.194087342373
			11'd198: out = 32'b00000000000000000001100011111000; // input=0.19384765625, output=0.195082689101
			11'd199: out = 32'b00000000000000000001100100011001; // input=0.19482421875, output=0.19607823163
			11'd200: out = 32'b00000000000000000001100100111010; // input=0.19580078125, output=0.19707397106
			11'd201: out = 32'b00000000000000000001100101011010; // input=0.19677734375, output=0.198069908498
			11'd202: out = 32'b00000000000000000001100101111011; // input=0.19775390625, output=0.19906604505
			11'd203: out = 32'b00000000000000000001100110011100; // input=0.19873046875, output=0.200062381825
			11'd204: out = 32'b00000000000000000001100110111100; // input=0.19970703125, output=0.201058919932
			11'd205: out = 32'b00000000000000000001100111011101; // input=0.20068359375, output=0.202055660484
			11'd206: out = 32'b00000000000000000001100111111110; // input=0.20166015625, output=0.203052604596
			11'd207: out = 32'b00000000000000000001101000011110; // input=0.20263671875, output=0.204049753384
			11'd208: out = 32'b00000000000000000001101000111111; // input=0.20361328125, output=0.205047107966
			11'd209: out = 32'b00000000000000000001101001100000; // input=0.20458984375, output=0.206044669461
			11'd210: out = 32'b00000000000000000001101010000000; // input=0.20556640625, output=0.207042438993
			11'd211: out = 32'b00000000000000000001101010100001; // input=0.20654296875, output=0.208040417685
			11'd212: out = 32'b00000000000000000001101011000010; // input=0.20751953125, output=0.209038606664
			11'd213: out = 32'b00000000000000000001101011100010; // input=0.20849609375, output=0.210037007058
			11'd214: out = 32'b00000000000000000001101100000011; // input=0.20947265625, output=0.211035619996
			11'd215: out = 32'b00000000000000000001101100100100; // input=0.21044921875, output=0.212034446612
			11'd216: out = 32'b00000000000000000001101101000101; // input=0.21142578125, output=0.21303348804
			11'd217: out = 32'b00000000000000000001101101100101; // input=0.21240234375, output=0.214032745416
			11'd218: out = 32'b00000000000000000001101110000110; // input=0.21337890625, output=0.215032219878
			11'd219: out = 32'b00000000000000000001101110100111; // input=0.21435546875, output=0.216031912567
			11'd220: out = 32'b00000000000000000001101111001000; // input=0.21533203125, output=0.217031824626
			11'd221: out = 32'b00000000000000000001101111101000; // input=0.21630859375, output=0.218031957201
			11'd222: out = 32'b00000000000000000001110000001001; // input=0.21728515625, output=0.219032311437
			11'd223: out = 32'b00000000000000000001110000101010; // input=0.21826171875, output=0.220032888484
			11'd224: out = 32'b00000000000000000001110001001011; // input=0.21923828125, output=0.221033689493
			11'd225: out = 32'b00000000000000000001110001101100; // input=0.22021484375, output=0.222034715618
			11'd226: out = 32'b00000000000000000001110010001100; // input=0.22119140625, output=0.223035968015
			11'd227: out = 32'b00000000000000000001110010101101; // input=0.22216796875, output=0.224037447841
			11'd228: out = 32'b00000000000000000001110011001110; // input=0.22314453125, output=0.225039156258
			11'd229: out = 32'b00000000000000000001110011101111; // input=0.22412109375, output=0.226041094426
			11'd230: out = 32'b00000000000000000001110100010000; // input=0.22509765625, output=0.227043263512
			11'd231: out = 32'b00000000000000000001110100110001; // input=0.22607421875, output=0.228045664681
			11'd232: out = 32'b00000000000000000001110101010001; // input=0.22705078125, output=0.229048299103
			11'd233: out = 32'b00000000000000000001110101110010; // input=0.22802734375, output=0.23005116795
			11'd234: out = 32'b00000000000000000001110110010011; // input=0.22900390625, output=0.231054272395
			11'd235: out = 32'b00000000000000000001110110110100; // input=0.22998046875, output=0.232057613615
			11'd236: out = 32'b00000000000000000001110111010101; // input=0.23095703125, output=0.233061192788
			11'd237: out = 32'b00000000000000000001110111110110; // input=0.23193359375, output=0.234065011095
			11'd238: out = 32'b00000000000000000001111000010111; // input=0.23291015625, output=0.23506906972
			11'd239: out = 32'b00000000000000000001111000111000; // input=0.23388671875, output=0.236073369847
			11'd240: out = 32'b00000000000000000001111001011001; // input=0.23486328125, output=0.237077912665
			11'd241: out = 32'b00000000000000000001111001111001; // input=0.23583984375, output=0.238082699365
			11'd242: out = 32'b00000000000000000001111010011010; // input=0.23681640625, output=0.239087731139
			11'd243: out = 32'b00000000000000000001111010111011; // input=0.23779296875, output=0.240093009183
			11'd244: out = 32'b00000000000000000001111011011100; // input=0.23876953125, output=0.241098534694
			11'd245: out = 32'b00000000000000000001111011111101; // input=0.23974609375, output=0.242104308872
			11'd246: out = 32'b00000000000000000001111100011110; // input=0.24072265625, output=0.243110332922
			11'd247: out = 32'b00000000000000000001111100111111; // input=0.24169921875, output=0.244116608046
			11'd248: out = 32'b00000000000000000001111101100000; // input=0.24267578125, output=0.245123135455
			11'd249: out = 32'b00000000000000000001111110000001; // input=0.24365234375, output=0.246129916357
			11'd250: out = 32'b00000000000000000001111110100010; // input=0.24462890625, output=0.247136951966
			11'd251: out = 32'b00000000000000000001111111000011; // input=0.24560546875, output=0.248144243497
			11'd252: out = 32'b00000000000000000001111111100100; // input=0.24658203125, output=0.249151792168
			11'd253: out = 32'b00000000000000000010000000000101; // input=0.24755859375, output=0.2501595992
			11'd254: out = 32'b00000000000000000010000000100110; // input=0.24853515625, output=0.251167665816
			11'd255: out = 32'b00000000000000000010000001000111; // input=0.24951171875, output=0.252175993242
			11'd256: out = 32'b00000000000000000010000001101000; // input=0.25048828125, output=0.253184582706
			11'd257: out = 32'b00000000000000000010000010001001; // input=0.25146484375, output=0.25419343544
			11'd258: out = 32'b00000000000000000010000010101010; // input=0.25244140625, output=0.255202552678
			11'd259: out = 32'b00000000000000000010000011001100; // input=0.25341796875, output=0.256211935655
			11'd260: out = 32'b00000000000000000010000011101101; // input=0.25439453125, output=0.257221585612
			11'd261: out = 32'b00000000000000000010000100001110; // input=0.25537109375, output=0.25823150379
			11'd262: out = 32'b00000000000000000010000100101111; // input=0.25634765625, output=0.259241691435
			11'd263: out = 32'b00000000000000000010000101010000; // input=0.25732421875, output=0.260252149793
			11'd264: out = 32'b00000000000000000010000101110001; // input=0.25830078125, output=0.261262880115
			11'd265: out = 32'b00000000000000000010000110010010; // input=0.25927734375, output=0.262273883654
			11'd266: out = 32'b00000000000000000010000110110011; // input=0.26025390625, output=0.263285161666
			11'd267: out = 32'b00000000000000000010000111010100; // input=0.26123046875, output=0.26429671541
			11'd268: out = 32'b00000000000000000010000111110110; // input=0.26220703125, output=0.265308546147
			11'd269: out = 32'b00000000000000000010001000010111; // input=0.26318359375, output=0.266320655141
			11'd270: out = 32'b00000000000000000010001000111000; // input=0.26416015625, output=0.267333043661
			11'd271: out = 32'b00000000000000000010001001011001; // input=0.26513671875, output=0.268345712975
			11'd272: out = 32'b00000000000000000010001001111010; // input=0.26611328125, output=0.269358664358
			11'd273: out = 32'b00000000000000000010001010011100; // input=0.26708984375, output=0.270371899086
			11'd274: out = 32'b00000000000000000010001010111101; // input=0.26806640625, output=0.271385418436
			11'd275: out = 32'b00000000000000000010001011011110; // input=0.26904296875, output=0.272399223693
			11'd276: out = 32'b00000000000000000010001011111111; // input=0.27001953125, output=0.273413316139
			11'd277: out = 32'b00000000000000000010001100100000; // input=0.27099609375, output=0.274427697064
			11'd278: out = 32'b00000000000000000010001101000010; // input=0.27197265625, output=0.275442367758
			11'd279: out = 32'b00000000000000000010001101100011; // input=0.27294921875, output=0.276457329516
			11'd280: out = 32'b00000000000000000010001110000100; // input=0.27392578125, output=0.277472583634
			11'd281: out = 32'b00000000000000000010001110100101; // input=0.27490234375, output=0.278488131412
			11'd282: out = 32'b00000000000000000010001111000111; // input=0.27587890625, output=0.279503974155
			11'd283: out = 32'b00000000000000000010001111101000; // input=0.27685546875, output=0.280520113167
			11'd284: out = 32'b00000000000000000010010000001001; // input=0.27783203125, output=0.28153654976
			11'd285: out = 32'b00000000000000000010010000101011; // input=0.27880859375, output=0.282553285244
			11'd286: out = 32'b00000000000000000010010001001100; // input=0.27978515625, output=0.283570320937
			11'd287: out = 32'b00000000000000000010010001101101; // input=0.28076171875, output=0.284587658157
			11'd288: out = 32'b00000000000000000010010010001111; // input=0.28173828125, output=0.285605298226
			11'd289: out = 32'b00000000000000000010010010110000; // input=0.28271484375, output=0.28662324247
			11'd290: out = 32'b00000000000000000010010011010001; // input=0.28369140625, output=0.287641492218
			11'd291: out = 32'b00000000000000000010010011110011; // input=0.28466796875, output=0.288660048801
			11'd292: out = 32'b00000000000000000010010100010100; // input=0.28564453125, output=0.289678913555
			11'd293: out = 32'b00000000000000000010010100110110; // input=0.28662109375, output=0.290698087817
			11'd294: out = 32'b00000000000000000010010101010111; // input=0.28759765625, output=0.291717572931
			11'd295: out = 32'b00000000000000000010010101111000; // input=0.28857421875, output=0.292737370241
			11'd296: out = 32'b00000000000000000010010110011010; // input=0.28955078125, output=0.293757481095
			11'd297: out = 32'b00000000000000000010010110111011; // input=0.29052734375, output=0.294777906847
			11'd298: out = 32'b00000000000000000010010111011101; // input=0.29150390625, output=0.29579864885
			11'd299: out = 32'b00000000000000000010010111111110; // input=0.29248046875, output=0.296819708463
			11'd300: out = 32'b00000000000000000010011000100000; // input=0.29345703125, output=0.29784108705
			11'd301: out = 32'b00000000000000000010011001000001; // input=0.29443359375, output=0.298862785975
			11'd302: out = 32'b00000000000000000010011001100011; // input=0.29541015625, output=0.299884806608
			11'd303: out = 32'b00000000000000000010011010000100; // input=0.29638671875, output=0.300907150321
			11'd304: out = 32'b00000000000000000010011010100110; // input=0.29736328125, output=0.30192981849
			11'd305: out = 32'b00000000000000000010011011000111; // input=0.29833984375, output=0.302952812495
			11'd306: out = 32'b00000000000000000010011011101001; // input=0.29931640625, output=0.30397613372
			11'd307: out = 32'b00000000000000000010011100001010; // input=0.30029296875, output=0.304999783551
			11'd308: out = 32'b00000000000000000010011100101100; // input=0.30126953125, output=0.306023763378
			11'd309: out = 32'b00000000000000000010011101001101; // input=0.30224609375, output=0.307048074597
			11'd310: out = 32'b00000000000000000010011101101111; // input=0.30322265625, output=0.308072718603
			11'd311: out = 32'b00000000000000000010011110010001; // input=0.30419921875, output=0.309097696799
			11'd312: out = 32'b00000000000000000010011110110010; // input=0.30517578125, output=0.310123010591
			11'd313: out = 32'b00000000000000000010011111010100; // input=0.30615234375, output=0.311148661385
			11'd314: out = 32'b00000000000000000010011111110101; // input=0.30712890625, output=0.312174650596
			11'd315: out = 32'b00000000000000000010100000010111; // input=0.30810546875, output=0.31320097964
			11'd316: out = 32'b00000000000000000010100000111001; // input=0.30908203125, output=0.314227649936
			11'd317: out = 32'b00000000000000000010100001011010; // input=0.31005859375, output=0.315254662909
			11'd318: out = 32'b00000000000000000010100001111100; // input=0.31103515625, output=0.316282019985
			11'd319: out = 32'b00000000000000000010100010011110; // input=0.31201171875, output=0.317309722597
			11'd320: out = 32'b00000000000000000010100010111111; // input=0.31298828125, output=0.318337772181
			11'd321: out = 32'b00000000000000000010100011100001; // input=0.31396484375, output=0.319366170175
			11'd322: out = 32'b00000000000000000010100100000011; // input=0.31494140625, output=0.320394918022
			11'd323: out = 32'b00000000000000000010100100100100; // input=0.31591796875, output=0.32142401717
			11'd324: out = 32'b00000000000000000010100101000110; // input=0.31689453125, output=0.32245346907
			11'd325: out = 32'b00000000000000000010100101101000; // input=0.31787109375, output=0.323483275177
			11'd326: out = 32'b00000000000000000010100110001010; // input=0.31884765625, output=0.32451343695
			11'd327: out = 32'b00000000000000000010100110101011; // input=0.31982421875, output=0.325543955852
			11'd328: out = 32'b00000000000000000010100111001101; // input=0.32080078125, output=0.326574833351
			11'd329: out = 32'b00000000000000000010100111101111; // input=0.32177734375, output=0.327606070917
			11'd330: out = 32'b00000000000000000010101000010001; // input=0.32275390625, output=0.328637670026
			11'd331: out = 32'b00000000000000000010101000110011; // input=0.32373046875, output=0.329669632158
			11'd332: out = 32'b00000000000000000010101001010100; // input=0.32470703125, output=0.330701958797
			11'd333: out = 32'b00000000000000000010101001110110; // input=0.32568359375, output=0.331734651429
			11'd334: out = 32'b00000000000000000010101010011000; // input=0.32666015625, output=0.332767711548
			11'd335: out = 32'b00000000000000000010101010111010; // input=0.32763671875, output=0.333801140649
			11'd336: out = 32'b00000000000000000010101011011100; // input=0.32861328125, output=0.334834940233
			11'd337: out = 32'b00000000000000000010101011111110; // input=0.32958984375, output=0.335869111804
			11'd338: out = 32'b00000000000000000010101100100000; // input=0.33056640625, output=0.336903656873
			11'd339: out = 32'b00000000000000000010101101000010; // input=0.33154296875, output=0.337938576951
			11'd340: out = 32'b00000000000000000010101101100011; // input=0.33251953125, output=0.338973873558
			11'd341: out = 32'b00000000000000000010101110000101; // input=0.33349609375, output=0.340009548215
			11'd342: out = 32'b00000000000000000010101110100111; // input=0.33447265625, output=0.341045602449
			11'd343: out = 32'b00000000000000000010101111001001; // input=0.33544921875, output=0.34208203779
			11'd344: out = 32'b00000000000000000010101111101011; // input=0.33642578125, output=0.343118855775
			11'd345: out = 32'b00000000000000000010110000001101; // input=0.33740234375, output=0.344156057942
			11'd346: out = 32'b00000000000000000010110000101111; // input=0.33837890625, output=0.345193645838
			11'd347: out = 32'b00000000000000000010110001010001; // input=0.33935546875, output=0.346231621009
			11'd348: out = 32'b00000000000000000010110001110011; // input=0.34033203125, output=0.347269985011
			11'd349: out = 32'b00000000000000000010110010010101; // input=0.34130859375, output=0.348308739401
			11'd350: out = 32'b00000000000000000010110010110111; // input=0.34228515625, output=0.349347885742
			11'd351: out = 32'b00000000000000000010110011011001; // input=0.34326171875, output=0.350387425601
			11'd352: out = 32'b00000000000000000010110011111100; // input=0.34423828125, output=0.351427360551
			11'd353: out = 32'b00000000000000000010110100011110; // input=0.34521484375, output=0.352467692167
			11'd354: out = 32'b00000000000000000010110101000000; // input=0.34619140625, output=0.353508422032
			11'd355: out = 32'b00000000000000000010110101100010; // input=0.34716796875, output=0.354549551733
			11'd356: out = 32'b00000000000000000010110110000100; // input=0.34814453125, output=0.355591082858
			11'd357: out = 32'b00000000000000000010110110100110; // input=0.34912109375, output=0.356633017006
			11'd358: out = 32'b00000000000000000010110111001000; // input=0.35009765625, output=0.357675355776
			11'd359: out = 32'b00000000000000000010110111101010; // input=0.35107421875, output=0.358718100774
			11'd360: out = 32'b00000000000000000010111000001101; // input=0.35205078125, output=0.359761253611
			11'd361: out = 32'b00000000000000000010111000101111; // input=0.35302734375, output=0.360804815901
			11'd362: out = 32'b00000000000000000010111001010001; // input=0.35400390625, output=0.361848789265
			11'd363: out = 32'b00000000000000000010111001110011; // input=0.35498046875, output=0.362893175329
			11'd364: out = 32'b00000000000000000010111010010110; // input=0.35595703125, output=0.363937975722
			11'd365: out = 32'b00000000000000000010111010111000; // input=0.35693359375, output=0.364983192081
			11'd366: out = 32'b00000000000000000010111011011010; // input=0.35791015625, output=0.366028826045
			11'd367: out = 32'b00000000000000000010111011111100; // input=0.35888671875, output=0.367074879261
			11'd368: out = 32'b00000000000000000010111100011111; // input=0.35986328125, output=0.368121353378
			11'd369: out = 32'b00000000000000000010111101000001; // input=0.36083984375, output=0.369168250053
			11'd370: out = 32'b00000000000000000010111101100011; // input=0.36181640625, output=0.370215570947
			11'd371: out = 32'b00000000000000000010111110000110; // input=0.36279296875, output=0.371263317726
			11'd372: out = 32'b00000000000000000010111110101000; // input=0.36376953125, output=0.372311492062
			11'd373: out = 32'b00000000000000000010111111001010; // input=0.36474609375, output=0.373360095631
			11'd374: out = 32'b00000000000000000010111111101101; // input=0.36572265625, output=0.374409130116
			11'd375: out = 32'b00000000000000000011000000001111; // input=0.36669921875, output=0.375458597205
			11'd376: out = 32'b00000000000000000011000000110001; // input=0.36767578125, output=0.37650849859
			11'd377: out = 32'b00000000000000000011000001010100; // input=0.36865234375, output=0.377558835969
			11'd378: out = 32'b00000000000000000011000001110110; // input=0.36962890625, output=0.378609611047
			11'd379: out = 32'b00000000000000000011000010011001; // input=0.37060546875, output=0.379660825532
			11'd380: out = 32'b00000000000000000011000010111011; // input=0.37158203125, output=0.38071248114
			11'd381: out = 32'b00000000000000000011000011011110; // input=0.37255859375, output=0.381764579591
			11'd382: out = 32'b00000000000000000011000100000000; // input=0.37353515625, output=0.38281712261
			11'd383: out = 32'b00000000000000000011000100100011; // input=0.37451171875, output=0.38387011193
			11'd384: out = 32'b00000000000000000011000101000101; // input=0.37548828125, output=0.384923549288
			11'd385: out = 32'b00000000000000000011000101101000; // input=0.37646484375, output=0.385977436426
			11'd386: out = 32'b00000000000000000011000110001010; // input=0.37744140625, output=0.387031775094
			11'd387: out = 32'b00000000000000000011000110101101; // input=0.37841796875, output=0.388086567045
			11'd388: out = 32'b00000000000000000011000111001111; // input=0.37939453125, output=0.38914181404
			11'd389: out = 32'b00000000000000000011000111110010; // input=0.38037109375, output=0.390197517845
			11'd390: out = 32'b00000000000000000011001000010101; // input=0.38134765625, output=0.391253680232
			11'd391: out = 32'b00000000000000000011001000110111; // input=0.38232421875, output=0.392310302978
			11'd392: out = 32'b00000000000000000011001001011010; // input=0.38330078125, output=0.393367387867
			11'd393: out = 32'b00000000000000000011001001111101; // input=0.38427734375, output=0.394424936689
			11'd394: out = 32'b00000000000000000011001010011111; // input=0.38525390625, output=0.395482951241
			11'd395: out = 32'b00000000000000000011001011000010; // input=0.38623046875, output=0.396541433322
			11'd396: out = 32'b00000000000000000011001011100101; // input=0.38720703125, output=0.397600384742
			11'd397: out = 32'b00000000000000000011001100000111; // input=0.38818359375, output=0.398659807314
			11'd398: out = 32'b00000000000000000011001100101010; // input=0.38916015625, output=0.399719702858
			11'd399: out = 32'b00000000000000000011001101001101; // input=0.39013671875, output=0.400780073201
			11'd400: out = 32'b00000000000000000011001101110000; // input=0.39111328125, output=0.401840920174
			11'd401: out = 32'b00000000000000000011001110010010; // input=0.39208984375, output=0.402902245618
			11'd402: out = 32'b00000000000000000011001110110101; // input=0.39306640625, output=0.403964051377
			11'd403: out = 32'b00000000000000000011001111011000; // input=0.39404296875, output=0.405026339302
			11'd404: out = 32'b00000000000000000011001111111011; // input=0.39501953125, output=0.406089111252
			11'd405: out = 32'b00000000000000000011010000011110; // input=0.39599609375, output=0.40715236909
			11'd406: out = 32'b00000000000000000011010001000000; // input=0.39697265625, output=0.408216114687
			11'd407: out = 32'b00000000000000000011010001100011; // input=0.39794921875, output=0.409280349921
			11'd408: out = 32'b00000000000000000011010010000110; // input=0.39892578125, output=0.410345076676
			11'd409: out = 32'b00000000000000000011010010101001; // input=0.39990234375, output=0.41141029684
			11'd410: out = 32'b00000000000000000011010011001100; // input=0.40087890625, output=0.412476012313
			11'd411: out = 32'b00000000000000000011010011101111; // input=0.40185546875, output=0.413542224997
			11'd412: out = 32'b00000000000000000011010100010010; // input=0.40283203125, output=0.414608936802
			11'd413: out = 32'b00000000000000000011010100110101; // input=0.40380859375, output=0.415676149646
			11'd414: out = 32'b00000000000000000011010101011000; // input=0.40478515625, output=0.416743865453
			11'd415: out = 32'b00000000000000000011010101111011; // input=0.40576171875, output=0.417812086153
			11'd416: out = 32'b00000000000000000011010110011110; // input=0.40673828125, output=0.418880813684
			11'd417: out = 32'b00000000000000000011010111000001; // input=0.40771484375, output=0.419950049991
			11'd418: out = 32'b00000000000000000011010111100100; // input=0.40869140625, output=0.421019797024
			11'd419: out = 32'b00000000000000000011011000000111; // input=0.40966796875, output=0.422090056743
			11'd420: out = 32'b00000000000000000011011000101010; // input=0.41064453125, output=0.423160831114
			11'd421: out = 32'b00000000000000000011011001001101; // input=0.41162109375, output=0.424232122107
			11'd422: out = 32'b00000000000000000011011001110000; // input=0.41259765625, output=0.425303931704
			11'd423: out = 32'b00000000000000000011011010010011; // input=0.41357421875, output=0.426376261892
			11'd424: out = 32'b00000000000000000011011010110111; // input=0.41455078125, output=0.427449114664
			11'd425: out = 32'b00000000000000000011011011011010; // input=0.41552734375, output=0.428522492022
			11'd426: out = 32'b00000000000000000011011011111101; // input=0.41650390625, output=0.429596395974
			11'd427: out = 32'b00000000000000000011011100100000; // input=0.41748046875, output=0.430670828538
			11'd428: out = 32'b00000000000000000011011101000011; // input=0.41845703125, output=0.431745791736
			11'd429: out = 32'b00000000000000000011011101100111; // input=0.41943359375, output=0.432821287599
			11'd430: out = 32'b00000000000000000011011110001010; // input=0.42041015625, output=0.433897318166
			11'd431: out = 32'b00000000000000000011011110101101; // input=0.42138671875, output=0.434973885483
			11'd432: out = 32'b00000000000000000011011111010001; // input=0.42236328125, output=0.436050991604
			11'd433: out = 32'b00000000000000000011011111110100; // input=0.42333984375, output=0.437128638589
			11'd434: out = 32'b00000000000000000011100000010111; // input=0.42431640625, output=0.438206828509
			11'd435: out = 32'b00000000000000000011100000111011; // input=0.42529296875, output=0.439285563439
			11'd436: out = 32'b00000000000000000011100001011110; // input=0.42626953125, output=0.440364845464
			11'd437: out = 32'b00000000000000000011100010000001; // input=0.42724609375, output=0.441444676676
			11'd438: out = 32'b00000000000000000011100010100101; // input=0.42822265625, output=0.442525059177
			11'd439: out = 32'b00000000000000000011100011001000; // input=0.42919921875, output=0.443605995073
			11'd440: out = 32'b00000000000000000011100011101100; // input=0.43017578125, output=0.444687486481
			11'd441: out = 32'b00000000000000000011100100001111; // input=0.43115234375, output=0.445769535526
			11'd442: out = 32'b00000000000000000011100100110010; // input=0.43212890625, output=0.446852144339
			11'd443: out = 32'b00000000000000000011100101010110; // input=0.43310546875, output=0.447935315062
			11'd444: out = 32'b00000000000000000011100101111001; // input=0.43408203125, output=0.449019049842
			11'd445: out = 32'b00000000000000000011100110011101; // input=0.43505859375, output=0.450103350837
			11'd446: out = 32'b00000000000000000011100111000001; // input=0.43603515625, output=0.451188220212
			11'd447: out = 32'b00000000000000000011100111100100; // input=0.43701171875, output=0.452273660141
			11'd448: out = 32'b00000000000000000011101000001000; // input=0.43798828125, output=0.453359672806
			11'd449: out = 32'b00000000000000000011101000101011; // input=0.43896484375, output=0.454446260396
			11'd450: out = 32'b00000000000000000011101001001111; // input=0.43994140625, output=0.455533425112
			11'd451: out = 32'b00000000000000000011101001110011; // input=0.44091796875, output=0.456621169161
			11'd452: out = 32'b00000000000000000011101010010110; // input=0.44189453125, output=0.457709494758
			11'd453: out = 32'b00000000000000000011101010111010; // input=0.44287109375, output=0.458798404129
			11'd454: out = 32'b00000000000000000011101011011110; // input=0.44384765625, output=0.459887899507
			11'd455: out = 32'b00000000000000000011101100000001; // input=0.44482421875, output=0.460977983136
			11'd456: out = 32'b00000000000000000011101100100101; // input=0.44580078125, output=0.462068657266
			11'd457: out = 32'b00000000000000000011101101001001; // input=0.44677734375, output=0.463159924156
			11'd458: out = 32'b00000000000000000011101101101101; // input=0.44775390625, output=0.464251786078
			11'd459: out = 32'b00000000000000000011101110010000; // input=0.44873046875, output=0.465344245308
			11'd460: out = 32'b00000000000000000011101110110100; // input=0.44970703125, output=0.466437304135
			11'd461: out = 32'b00000000000000000011101111011000; // input=0.45068359375, output=0.467530964854
			11'd462: out = 32'b00000000000000000011101111111100; // input=0.45166015625, output=0.468625229772
			11'd463: out = 32'b00000000000000000011110000100000; // input=0.45263671875, output=0.469720101202
			11'd464: out = 32'b00000000000000000011110001000100; // input=0.45361328125, output=0.47081558147
			11'd465: out = 32'b00000000000000000011110001101000; // input=0.45458984375, output=0.47191167291
			11'd466: out = 32'b00000000000000000011110010001100; // input=0.45556640625, output=0.473008377863
			11'd467: out = 32'b00000000000000000011110010101111; // input=0.45654296875, output=0.474105698684
			11'd468: out = 32'b00000000000000000011110011010011; // input=0.45751953125, output=0.475203637734
			11'd469: out = 32'b00000000000000000011110011110111; // input=0.45849609375, output=0.476302197385
			11'd470: out = 32'b00000000000000000011110100011011; // input=0.45947265625, output=0.477401380019
			11'd471: out = 32'b00000000000000000011110101000000; // input=0.46044921875, output=0.478501188027
			11'd472: out = 32'b00000000000000000011110101100100; // input=0.46142578125, output=0.47960162381
			11'd473: out = 32'b00000000000000000011110110001000; // input=0.46240234375, output=0.48070268978
			11'd474: out = 32'b00000000000000000011110110101100; // input=0.46337890625, output=0.481804388357
			11'd475: out = 32'b00000000000000000011110111010000; // input=0.46435546875, output=0.482906721972
			11'd476: out = 32'b00000000000000000011110111110100; // input=0.46533203125, output=0.484009693068
			11'd477: out = 32'b00000000000000000011111000011000; // input=0.46630859375, output=0.485113304095
			11'd478: out = 32'b00000000000000000011111000111100; // input=0.46728515625, output=0.486217557514
			11'd479: out = 32'b00000000000000000011111001100001; // input=0.46826171875, output=0.487322455798
			11'd480: out = 32'b00000000000000000011111010000101; // input=0.46923828125, output=0.48842800143
			11'd481: out = 32'b00000000000000000011111010101001; // input=0.47021484375, output=0.489534196901
			11'd482: out = 32'b00000000000000000011111011001101; // input=0.47119140625, output=0.490641044716
			11'd483: out = 32'b00000000000000000011111011110010; // input=0.47216796875, output=0.491748547388
			11'd484: out = 32'b00000000000000000011111100010110; // input=0.47314453125, output=0.492856707441
			11'd485: out = 32'b00000000000000000011111100111010; // input=0.47412109375, output=0.493965527411
			11'd486: out = 32'b00000000000000000011111101011111; // input=0.47509765625, output=0.495075009844
			11'd487: out = 32'b00000000000000000011111110000011; // input=0.47607421875, output=0.496185157297
			11'd488: out = 32'b00000000000000000011111110100111; // input=0.47705078125, output=0.497295972337
			11'd489: out = 32'b00000000000000000011111111001100; // input=0.47802734375, output=0.498407457545
			11'd490: out = 32'b00000000000000000011111111110000; // input=0.47900390625, output=0.499519615509
			11'd491: out = 32'b00000000000000000100000000010101; // input=0.47998046875, output=0.500632448832
			11'd492: out = 32'b00000000000000000100000000111001; // input=0.48095703125, output=0.501745960124
			11'd493: out = 32'b00000000000000000100000001011110; // input=0.48193359375, output=0.502860152012
			11'd494: out = 32'b00000000000000000100000010000010; // input=0.48291015625, output=0.503975027128
			11'd495: out = 32'b00000000000000000100000010100111; // input=0.48388671875, output=0.505090588121
			11'd496: out = 32'b00000000000000000100000011001011; // input=0.48486328125, output=0.506206837649
			11'd497: out = 32'b00000000000000000100000011110000; // input=0.48583984375, output=0.50732377838
			11'd498: out = 32'b00000000000000000100000100010101; // input=0.48681640625, output=0.508441412998
			11'd499: out = 32'b00000000000000000100000100111001; // input=0.48779296875, output=0.509559744196
			11'd500: out = 32'b00000000000000000100000101011110; // input=0.48876953125, output=0.510678774679
			11'd501: out = 32'b00000000000000000100000110000011; // input=0.48974609375, output=0.511798507164
			11'd502: out = 32'b00000000000000000100000110100111; // input=0.49072265625, output=0.51291894438
			11'd503: out = 32'b00000000000000000100000111001100; // input=0.49169921875, output=0.51404008907
			11'd504: out = 32'b00000000000000000100000111110001; // input=0.49267578125, output=0.515161943987
			11'd505: out = 32'b00000000000000000100001000010110; // input=0.49365234375, output=0.516284511897
			11'd506: out = 32'b00000000000000000100001000111010; // input=0.49462890625, output=0.517407795578
			11'd507: out = 32'b00000000000000000100001001011111; // input=0.49560546875, output=0.518531797822
			11'd508: out = 32'b00000000000000000100001010000100; // input=0.49658203125, output=0.519656521432
			11'd509: out = 32'b00000000000000000100001010101001; // input=0.49755859375, output=0.520781969224
			11'd510: out = 32'b00000000000000000100001011001110; // input=0.49853515625, output=0.521908144027
			11'd511: out = 32'b00000000000000000100001011110011; // input=0.49951171875, output=0.523035048684
			11'd512: out = 32'b00000000000000000100001100011000; // input=0.50048828125, output=0.524162686048
			11'd513: out = 32'b00000000000000000100001100111101; // input=0.50146484375, output=0.525291058987
			11'd514: out = 32'b00000000000000000100001101100010; // input=0.50244140625, output=0.526420170383
			11'd515: out = 32'b00000000000000000100001110000111; // input=0.50341796875, output=0.527550023129
			11'd516: out = 32'b00000000000000000100001110101100; // input=0.50439453125, output=0.528680620133
			11'd517: out = 32'b00000000000000000100001111010001; // input=0.50537109375, output=0.529811964315
			11'd518: out = 32'b00000000000000000100001111110110; // input=0.50634765625, output=0.53094405861
			11'd519: out = 32'b00000000000000000100010000011011; // input=0.50732421875, output=0.532076905965
			11'd520: out = 32'b00000000000000000100010001000000; // input=0.50830078125, output=0.533210509343
			11'd521: out = 32'b00000000000000000100010001100101; // input=0.50927734375, output=0.534344871718
			11'd522: out = 32'b00000000000000000100010010001011; // input=0.51025390625, output=0.53547999608
			11'd523: out = 32'b00000000000000000100010010110000; // input=0.51123046875, output=0.536615885432
			11'd524: out = 32'b00000000000000000100010011010101; // input=0.51220703125, output=0.537752542791
			11'd525: out = 32'b00000000000000000100010011111010; // input=0.51318359375, output=0.538889971188
			11'd526: out = 32'b00000000000000000100010100100000; // input=0.51416015625, output=0.54002817367
			11'd527: out = 32'b00000000000000000100010101000101; // input=0.51513671875, output=0.541167153296
			11'd528: out = 32'b00000000000000000100010101101010; // input=0.51611328125, output=0.542306913141
			11'd529: out = 32'b00000000000000000100010110010000; // input=0.51708984375, output=0.543447456295
			11'd530: out = 32'b00000000000000000100010110110101; // input=0.51806640625, output=0.544588785861
			11'd531: out = 32'b00000000000000000100010111011011; // input=0.51904296875, output=0.545730904958
			11'd532: out = 32'b00000000000000000100011000000000; // input=0.52001953125, output=0.54687381672
			11'd533: out = 32'b00000000000000000100011000100101; // input=0.52099609375, output=0.548017524295
			11'd534: out = 32'b00000000000000000100011001001011; // input=0.52197265625, output=0.549162030848
			11'd535: out = 32'b00000000000000000100011001110000; // input=0.52294921875, output=0.550307339557
			11'd536: out = 32'b00000000000000000100011010010110; // input=0.52392578125, output=0.551453453618
			11'd537: out = 32'b00000000000000000100011010111100; // input=0.52490234375, output=0.55260037624
			11'd538: out = 32'b00000000000000000100011011100001; // input=0.52587890625, output=0.553748110648
			11'd539: out = 32'b00000000000000000100011100000111; // input=0.52685546875, output=0.554896660084
			11'd540: out = 32'b00000000000000000100011100101101; // input=0.52783203125, output=0.556046027806
			11'd541: out = 32'b00000000000000000100011101010010; // input=0.52880859375, output=0.557196217085
			11'd542: out = 32'b00000000000000000100011101111000; // input=0.52978515625, output=0.558347231212
			11'd543: out = 32'b00000000000000000100011110011110; // input=0.53076171875, output=0.559499073492
			11'd544: out = 32'b00000000000000000100011111000011; // input=0.53173828125, output=0.560651747246
			11'd545: out = 32'b00000000000000000100011111101001; // input=0.53271484375, output=0.561805255813
			11'd546: out = 32'b00000000000000000100100000001111; // input=0.53369140625, output=0.562959602546
			11'd547: out = 32'b00000000000000000100100000110101; // input=0.53466796875, output=0.564114790818
			11'd548: out = 32'b00000000000000000100100001011011; // input=0.53564453125, output=0.565270824016
			11'd549: out = 32'b00000000000000000100100010000001; // input=0.53662109375, output=0.566427705546
			11'd550: out = 32'b00000000000000000100100010100111; // input=0.53759765625, output=0.567585438829
			11'd551: out = 32'b00000000000000000100100011001101; // input=0.53857421875, output=0.568744027306
			11'd552: out = 32'b00000000000000000100100011110011; // input=0.53955078125, output=0.569903474432
			11'd553: out = 32'b00000000000000000100100100011001; // input=0.54052734375, output=0.571063783681
			11'd554: out = 32'b00000000000000000100100100111111; // input=0.54150390625, output=0.572224958546
			11'd555: out = 32'b00000000000000000100100101100101; // input=0.54248046875, output=0.573387002535
			11'd556: out = 32'b00000000000000000100100110001011; // input=0.54345703125, output=0.574549919176
			11'd557: out = 32'b00000000000000000100100110110001; // input=0.54443359375, output=0.575713712013
			11'd558: out = 32'b00000000000000000100100111010111; // input=0.54541015625, output=0.576878384612
			11'd559: out = 32'b00000000000000000100100111111101; // input=0.54638671875, output=0.578043940552
			11'd560: out = 32'b00000000000000000100101000100100; // input=0.54736328125, output=0.579210383434
			11'd561: out = 32'b00000000000000000100101001001010; // input=0.54833984375, output=0.580377716876
			11'd562: out = 32'b00000000000000000100101001110000; // input=0.54931640625, output=0.581545944516
			11'd563: out = 32'b00000000000000000100101010010110; // input=0.55029296875, output=0.58271507001
			11'd564: out = 32'b00000000000000000100101010111101; // input=0.55126953125, output=0.583885097033
			11'd565: out = 32'b00000000000000000100101011100011; // input=0.55224609375, output=0.585056029278
			11'd566: out = 32'b00000000000000000100101100001010; // input=0.55322265625, output=0.586227870461
			11'd567: out = 32'b00000000000000000100101100110000; // input=0.55419921875, output=0.587400624313
			11'd568: out = 32'b00000000000000000100101101010110; // input=0.55517578125, output=0.588574294586
			11'd569: out = 32'b00000000000000000100101101111101; // input=0.55615234375, output=0.589748885055
			11'd570: out = 32'b00000000000000000100101110100011; // input=0.55712890625, output=0.590924399509
			11'd571: out = 32'b00000000000000000100101111001010; // input=0.55810546875, output=0.592100841762
			11'd572: out = 32'b00000000000000000100101111110001; // input=0.55908203125, output=0.593278215646
			11'd573: out = 32'b00000000000000000100110000010111; // input=0.56005859375, output=0.594456525014
			11'd574: out = 32'b00000000000000000100110000111110; // input=0.56103515625, output=0.595635773739
			11'd575: out = 32'b00000000000000000100110001100100; // input=0.56201171875, output=0.596815965716
			11'd576: out = 32'b00000000000000000100110010001011; // input=0.56298828125, output=0.597997104858
			11'd577: out = 32'b00000000000000000100110010110010; // input=0.56396484375, output=0.599179195102
			11'd578: out = 32'b00000000000000000100110011011001; // input=0.56494140625, output=0.600362240405
			11'd579: out = 32'b00000000000000000100110011111111; // input=0.56591796875, output=0.601546244745
			11'd580: out = 32'b00000000000000000100110100100110; // input=0.56689453125, output=0.602731212123
			11'd581: out = 32'b00000000000000000100110101001101; // input=0.56787109375, output=0.60391714656
			11'd582: out = 32'b00000000000000000100110101110100; // input=0.56884765625, output=0.6051040521
			11'd583: out = 32'b00000000000000000100110110011011; // input=0.56982421875, output=0.606291932808
			11'd584: out = 32'b00000000000000000100110111000010; // input=0.57080078125, output=0.607480792772
			11'd585: out = 32'b00000000000000000100110111101001; // input=0.57177734375, output=0.608670636103
			11'd586: out = 32'b00000000000000000100111000010000; // input=0.57275390625, output=0.609861466933
			11'd587: out = 32'b00000000000000000100111000110111; // input=0.57373046875, output=0.611053289418
			11'd588: out = 32'b00000000000000000100111001011110; // input=0.57470703125, output=0.612246107738
			11'd589: out = 32'b00000000000000000100111010000101; // input=0.57568359375, output=0.613439926093
			11'd590: out = 32'b00000000000000000100111010101100; // input=0.57666015625, output=0.614634748708
			11'd591: out = 32'b00000000000000000100111011010100; // input=0.57763671875, output=0.615830579834
			11'd592: out = 32'b00000000000000000100111011111011; // input=0.57861328125, output=0.617027423741
			11'd593: out = 32'b00000000000000000100111100100010; // input=0.57958984375, output=0.618225284727
			11'd594: out = 32'b00000000000000000100111101001001; // input=0.58056640625, output=0.619424167112
			11'd595: out = 32'b00000000000000000100111101110001; // input=0.58154296875, output=0.62062407524
			11'd596: out = 32'b00000000000000000100111110011000; // input=0.58251953125, output=0.621825013482
			11'd597: out = 32'b00000000000000000100111110111111; // input=0.58349609375, output=0.623026986232
			11'd598: out = 32'b00000000000000000100111111100111; // input=0.58447265625, output=0.624229997907
			11'd599: out = 32'b00000000000000000101000000001110; // input=0.58544921875, output=0.625434052954
			11'd600: out = 32'b00000000000000000101000000110110; // input=0.58642578125, output=0.62663915584
			11'd601: out = 32'b00000000000000000101000001011101; // input=0.58740234375, output=0.627845311062
			11'd602: out = 32'b00000000000000000101000010000101; // input=0.58837890625, output=0.629052523141
			11'd603: out = 32'b00000000000000000101000010101100; // input=0.58935546875, output=0.630260796623
			11'd604: out = 32'b00000000000000000101000011010100; // input=0.59033203125, output=0.631470136082
			11'd605: out = 32'b00000000000000000101000011111100; // input=0.59130859375, output=0.632680546116
			11'd606: out = 32'b00000000000000000101000100100011; // input=0.59228515625, output=0.633892031354
			11'd607: out = 32'b00000000000000000101000101001011; // input=0.59326171875, output=0.635104596447
			11'd608: out = 32'b00000000000000000101000101110011; // input=0.59423828125, output=0.636318246077
			11'd609: out = 32'b00000000000000000101000110011011; // input=0.59521484375, output=0.63753298495
			11'd610: out = 32'b00000000000000000101000111000011; // input=0.59619140625, output=0.638748817803
			11'd611: out = 32'b00000000000000000101000111101010; // input=0.59716796875, output=0.639965749399
			11'd612: out = 32'b00000000000000000101001000010010; // input=0.59814453125, output=0.641183784528
			11'd613: out = 32'b00000000000000000101001000111010; // input=0.59912109375, output=0.64240292801
			11'd614: out = 32'b00000000000000000101001001100010; // input=0.60009765625, output=0.643623184695
			11'd615: out = 32'b00000000000000000101001010001010; // input=0.60107421875, output=0.644844559457
			11'd616: out = 32'b00000000000000000101001010110010; // input=0.60205078125, output=0.646067057204
			11'd617: out = 32'b00000000000000000101001011011010; // input=0.60302734375, output=0.647290682871
			11'd618: out = 32'b00000000000000000101001100000011; // input=0.60400390625, output=0.648515441423
			11'd619: out = 32'b00000000000000000101001100101011; // input=0.60498046875, output=0.649741337855
			11'd620: out = 32'b00000000000000000101001101010011; // input=0.60595703125, output=0.650968377191
			11'd621: out = 32'b00000000000000000101001101111011; // input=0.60693359375, output=0.652196564486
			11'd622: out = 32'b00000000000000000101001110100011; // input=0.60791015625, output=0.653425904828
			11'd623: out = 32'b00000000000000000101001111001100; // input=0.60888671875, output=0.654656403331
			11'd624: out = 32'b00000000000000000101001111110100; // input=0.60986328125, output=0.655888065144
			11'd625: out = 32'b00000000000000000101010000011101; // input=0.61083984375, output=0.657120895447
			11'd626: out = 32'b00000000000000000101010001000101; // input=0.61181640625, output=0.658354899451
			11'd627: out = 32'b00000000000000000101010001101101; // input=0.61279296875, output=0.659590082398
			11'd628: out = 32'b00000000000000000101010010010110; // input=0.61376953125, output=0.660826449565
			11'd629: out = 32'b00000000000000000101010010111111; // input=0.61474609375, output=0.662064006259
			11'd630: out = 32'b00000000000000000101010011100111; // input=0.61572265625, output=0.66330275782
			11'd631: out = 32'b00000000000000000101010100010000; // input=0.61669921875, output=0.664542709624
			11'd632: out = 32'b00000000000000000101010100111000; // input=0.61767578125, output=0.665783867077
			11'd633: out = 32'b00000000000000000101010101100001; // input=0.61865234375, output=0.667026235621
			11'd634: out = 32'b00000000000000000101010110001010; // input=0.61962890625, output=0.668269820732
			11'd635: out = 32'b00000000000000000101010110110011; // input=0.62060546875, output=0.669514627918
			11'd636: out = 32'b00000000000000000101010111011011; // input=0.62158203125, output=0.670760662725
			11'd637: out = 32'b00000000000000000101011000000100; // input=0.62255859375, output=0.672007930733
			11'd638: out = 32'b00000000000000000101011000101101; // input=0.62353515625, output=0.673256437555
			11'd639: out = 32'b00000000000000000101011001010110; // input=0.62451171875, output=0.674506188843
			11'd640: out = 32'b00000000000000000101011001111111; // input=0.62548828125, output=0.675757190283
			11'd641: out = 32'b00000000000000000101011010101000; // input=0.62646484375, output=0.677009447598
			11'd642: out = 32'b00000000000000000101011011010001; // input=0.62744140625, output=0.678262966548
			11'd643: out = 32'b00000000000000000101011011111010; // input=0.62841796875, output=0.679517752929
			11'd644: out = 32'b00000000000000000101011100100100; // input=0.62939453125, output=0.680773812575
			11'd645: out = 32'b00000000000000000101011101001101; // input=0.63037109375, output=0.682031151358
			11'd646: out = 32'b00000000000000000101011101110110; // input=0.63134765625, output=0.683289775188
			11'd647: out = 32'b00000000000000000101011110011111; // input=0.63232421875, output=0.684549690012
			11'd648: out = 32'b00000000000000000101011111001001; // input=0.63330078125, output=0.685810901818
			11'd649: out = 32'b00000000000000000101011111110010; // input=0.63427734375, output=0.687073416632
			11'd650: out = 32'b00000000000000000101100000011011; // input=0.63525390625, output=0.688337240519
			11'd651: out = 32'b00000000000000000101100001000101; // input=0.63623046875, output=0.689602379584
			11'd652: out = 32'b00000000000000000101100001101110; // input=0.63720703125, output=0.690868839974
			11'd653: out = 32'b00000000000000000101100010011000; // input=0.63818359375, output=0.692136627875
			11'd654: out = 32'b00000000000000000101100011000010; // input=0.63916015625, output=0.693405749514
			11'd655: out = 32'b00000000000000000101100011101011; // input=0.64013671875, output=0.694676211161
			11'd656: out = 32'b00000000000000000101100100010101; // input=0.64111328125, output=0.695948019125
			11'd657: out = 32'b00000000000000000101100100111111; // input=0.64208984375, output=0.697221179759
			11'd658: out = 32'b00000000000000000101100101101000; // input=0.64306640625, output=0.69849569946
			11'd659: out = 32'b00000000000000000101100110010010; // input=0.64404296875, output=0.699771584666
			11'd660: out = 32'b00000000000000000101100110111100; // input=0.64501953125, output=0.701048841859
			11'd661: out = 32'b00000000000000000101100111100110; // input=0.64599609375, output=0.702327477564
			11'd662: out = 32'b00000000000000000101101000010000; // input=0.64697265625, output=0.703607498353
			11'd663: out = 32'b00000000000000000101101000111010; // input=0.64794921875, output=0.70488891084
			11'd664: out = 32'b00000000000000000101101001100100; // input=0.64892578125, output=0.706171721686
			11'd665: out = 32'b00000000000000000101101010001110; // input=0.64990234375, output=0.707455937596
			11'd666: out = 32'b00000000000000000101101010111000; // input=0.65087890625, output=0.708741565323
			11'd667: out = 32'b00000000000000000101101011100010; // input=0.65185546875, output=0.710028611664
			11'd668: out = 32'b00000000000000000101101100001100; // input=0.65283203125, output=0.711317083466
			11'd669: out = 32'b00000000000000000101101100110111; // input=0.65380859375, output=0.712606987621
			11'd670: out = 32'b00000000000000000101101101100001; // input=0.65478515625, output=0.713898331071
			11'd671: out = 32'b00000000000000000101101110001011; // input=0.65576171875, output=0.715191120804
			11'd672: out = 32'b00000000000000000101101110110110; // input=0.65673828125, output=0.71648536386
			11'd673: out = 32'b00000000000000000101101111100000; // input=0.65771484375, output=0.717781067325
			11'd674: out = 32'b00000000000000000101110000001011; // input=0.65869140625, output=0.719078238338
			11'd675: out = 32'b00000000000000000101110000110101; // input=0.65966796875, output=0.720376884086
			11'd676: out = 32'b00000000000000000101110001100000; // input=0.66064453125, output=0.721677011809
			11'd677: out = 32'b00000000000000000101110010001011; // input=0.66162109375, output=0.722978628796
			11'd678: out = 32'b00000000000000000101110010110101; // input=0.66259765625, output=0.72428174239
			11'd679: out = 32'b00000000000000000101110011100000; // input=0.66357421875, output=0.725586359986
			11'd680: out = 32'b00000000000000000101110100001011; // input=0.66455078125, output=0.726892489032
			11'd681: out = 32'b00000000000000000101110100110110; // input=0.66552734375, output=0.728200137029
			11'd682: out = 32'b00000000000000000101110101100001; // input=0.66650390625, output=0.729509311532
			11'd683: out = 32'b00000000000000000101110110001100; // input=0.66748046875, output=0.730820020153
			11'd684: out = 32'b00000000000000000101110110110111; // input=0.66845703125, output=0.732132270556
			11'd685: out = 32'b00000000000000000101110111100010; // input=0.66943359375, output=0.733446070462
			11'd686: out = 32'b00000000000000000101111000001101; // input=0.67041015625, output=0.734761427651
			11'd687: out = 32'b00000000000000000101111000111000; // input=0.67138671875, output=0.736078349955
			11'd688: out = 32'b00000000000000000101111001100011; // input=0.67236328125, output=0.737396845268
			11'd689: out = 32'b00000000000000000101111010001110; // input=0.67333984375, output=0.73871692154
			11'd690: out = 32'b00000000000000000101111010111010; // input=0.67431640625, output=0.74003858678
			11'd691: out = 32'b00000000000000000101111011100101; // input=0.67529296875, output=0.741361849058
			11'd692: out = 32'b00000000000000000101111100010000; // input=0.67626953125, output=0.742686716502
			11'd693: out = 32'b00000000000000000101111100111100; // input=0.67724609375, output=0.744013197301
			11'd694: out = 32'b00000000000000000101111101100111; // input=0.67822265625, output=0.745341299708
			11'd695: out = 32'b00000000000000000101111110010011; // input=0.67919921875, output=0.746671032034
			11'd696: out = 32'b00000000000000000101111110111111; // input=0.68017578125, output=0.748002402655
			11'd697: out = 32'b00000000000000000101111111101010; // input=0.68115234375, output=0.749335420011
			11'd698: out = 32'b00000000000000000110000000010110; // input=0.68212890625, output=0.750670092604
			11'd699: out = 32'b00000000000000000110000001000010; // input=0.68310546875, output=0.752006429003
			11'd700: out = 32'b00000000000000000110000001101110; // input=0.68408203125, output=0.75334443784
			11'd701: out = 32'b00000000000000000110000010011001; // input=0.68505859375, output=0.754684127815
			11'd702: out = 32'b00000000000000000110000011000101; // input=0.68603515625, output=0.756025507694
			11'd703: out = 32'b00000000000000000110000011110001; // input=0.68701171875, output=0.757368586311
			11'd704: out = 32'b00000000000000000110000100011110; // input=0.68798828125, output=0.758713372569
			11'd705: out = 32'b00000000000000000110000101001010; // input=0.68896484375, output=0.760059875439
			11'd706: out = 32'b00000000000000000110000101110110; // input=0.68994140625, output=0.761408103962
			11'd707: out = 32'b00000000000000000110000110100010; // input=0.69091796875, output=0.76275806725
			11'd708: out = 32'b00000000000000000110000111001110; // input=0.69189453125, output=0.764109774486
			11'd709: out = 32'b00000000000000000110000111111011; // input=0.69287109375, output=0.765463234926
			11'd710: out = 32'b00000000000000000110001000100111; // input=0.69384765625, output=0.766818457899
			11'd711: out = 32'b00000000000000000110001001010100; // input=0.69482421875, output=0.768175452807
			11'd712: out = 32'b00000000000000000110001010000000; // input=0.69580078125, output=0.769534229128
			11'd713: out = 32'b00000000000000000110001010101101; // input=0.69677734375, output=0.770894796414
			11'd714: out = 32'b00000000000000000110001011011001; // input=0.69775390625, output=0.772257164294
			11'd715: out = 32'b00000000000000000110001100000110; // input=0.69873046875, output=0.773621342475
			11'd716: out = 32'b00000000000000000110001100110011; // input=0.69970703125, output=0.774987340742
			11'd717: out = 32'b00000000000000000110001101100000; // input=0.70068359375, output=0.776355168958
			11'd718: out = 32'b00000000000000000110001110001100; // input=0.70166015625, output=0.777724837066
			11'd719: out = 32'b00000000000000000110001110111001; // input=0.70263671875, output=0.779096355093
			11'd720: out = 32'b00000000000000000110001111100110; // input=0.70361328125, output=0.780469733143
			11'd721: out = 32'b00000000000000000110010000010011; // input=0.70458984375, output=0.781844981407
			11'd722: out = 32'b00000000000000000110010001000001; // input=0.70556640625, output=0.783222110157
			11'd723: out = 32'b00000000000000000110010001101110; // input=0.70654296875, output=0.78460112975
			11'd724: out = 32'b00000000000000000110010010011011; // input=0.70751953125, output=0.78598205063
			11'd725: out = 32'b00000000000000000110010011001000; // input=0.70849609375, output=0.787364883328
			11'd726: out = 32'b00000000000000000110010011110110; // input=0.70947265625, output=0.788749638461
			11'd727: out = 32'b00000000000000000110010100100011; // input=0.71044921875, output=0.790136326735
			11'd728: out = 32'b00000000000000000110010101010001; // input=0.71142578125, output=0.791524958947
			11'd729: out = 32'b00000000000000000110010101111110; // input=0.71240234375, output=0.792915545985
			11'd730: out = 32'b00000000000000000110010110101100; // input=0.71337890625, output=0.794308098827
			11'd731: out = 32'b00000000000000000110010111011010; // input=0.71435546875, output=0.795702628547
			11'd732: out = 32'b00000000000000000110011000000111; // input=0.71533203125, output=0.797099146312
			11'd733: out = 32'b00000000000000000110011000110101; // input=0.71630859375, output=0.798497663382
			11'd734: out = 32'b00000000000000000110011001100011; // input=0.71728515625, output=0.799898191117
			11'd735: out = 32'b00000000000000000110011010010001; // input=0.71826171875, output=0.801300740973
			11'd736: out = 32'b00000000000000000110011010111111; // input=0.71923828125, output=0.802705324505
			11'd737: out = 32'b00000000000000000110011011101101; // input=0.72021484375, output=0.804111953369
			11'd738: out = 32'b00000000000000000110011100011011; // input=0.72119140625, output=0.805520639322
			11'd739: out = 32'b00000000000000000110011101001010; // input=0.72216796875, output=0.806931394221
			11'd740: out = 32'b00000000000000000110011101111000; // input=0.72314453125, output=0.808344230032
			11'd741: out = 32'b00000000000000000110011110100110; // input=0.72412109375, output=0.809759158821
			11'd742: out = 32'b00000000000000000110011111010101; // input=0.72509765625, output=0.811176192763
			11'd743: out = 32'b00000000000000000110100000000011; // input=0.72607421875, output=0.812595344141
			11'd744: out = 32'b00000000000000000110100000110010; // input=0.72705078125, output=0.814016625347
			11'd745: out = 32'b00000000000000000110100001100000; // input=0.72802734375, output=0.815440048882
			11'd746: out = 32'b00000000000000000110100010001111; // input=0.72900390625, output=0.816865627361
			11'd747: out = 32'b00000000000000000110100010111110; // input=0.72998046875, output=0.81829337351
			11'd748: out = 32'b00000000000000000110100011101101; // input=0.73095703125, output=0.819723300173
			11'd749: out = 32'b00000000000000000110100100011100; // input=0.73193359375, output=0.821155420307
			11'd750: out = 32'b00000000000000000110100101001011; // input=0.73291015625, output=0.822589746989
			11'd751: out = 32'b00000000000000000110100101111010; // input=0.73388671875, output=0.824026293413
			11'd752: out = 32'b00000000000000000110100110101001; // input=0.73486328125, output=0.825465072897
			11'd753: out = 32'b00000000000000000110100111011000; // input=0.73583984375, output=0.826906098877
			11'd754: out = 32'b00000000000000000110101000000111; // input=0.73681640625, output=0.828349384918
			11'd755: out = 32'b00000000000000000110101000110111; // input=0.73779296875, output=0.829794944707
			11'd756: out = 32'b00000000000000000110101001100110; // input=0.73876953125, output=0.831242792059
			11'd757: out = 32'b00000000000000000110101010010110; // input=0.73974609375, output=0.832692940918
			11'd758: out = 32'b00000000000000000110101011000101; // input=0.74072265625, output=0.834145405359
			11'd759: out = 32'b00000000000000000110101011110101; // input=0.74169921875, output=0.835600199588
			11'd760: out = 32'b00000000000000000110101100100101; // input=0.74267578125, output=0.837057337948
			11'd761: out = 32'b00000000000000000110101101010101; // input=0.74365234375, output=0.838516834915
			11'd762: out = 32'b00000000000000000110101110000100; // input=0.74462890625, output=0.839978705103
			11'd763: out = 32'b00000000000000000110101110110100; // input=0.74560546875, output=0.841442963267
			11'd764: out = 32'b00000000000000000110101111100100; // input=0.74658203125, output=0.842909624303
			11'd765: out = 32'b00000000000000000110110000010101; // input=0.74755859375, output=0.844378703249
			11'd766: out = 32'b00000000000000000110110001000101; // input=0.74853515625, output=0.845850215289
			11'd767: out = 32'b00000000000000000110110001110101; // input=0.74951171875, output=0.847324175756
			11'd768: out = 32'b00000000000000000110110010100101; // input=0.75048828125, output=0.84880060013
			11'd769: out = 32'b00000000000000000110110011010110; // input=0.75146484375, output=0.850279504044
			11'd770: out = 32'b00000000000000000110110100000111; // input=0.75244140625, output=0.851760903282
			11'd771: out = 32'b00000000000000000110110100110111; // input=0.75341796875, output=0.853244813787
			11'd772: out = 32'b00000000000000000110110101101000; // input=0.75439453125, output=0.854731251657
			11'd773: out = 32'b00000000000000000110110110011001; // input=0.75537109375, output=0.856220233152
			11'd774: out = 32'b00000000000000000110110111001001; // input=0.75634765625, output=0.857711774692
			11'd775: out = 32'b00000000000000000110110111111010; // input=0.75732421875, output=0.859205892863
			11'd776: out = 32'b00000000000000000110111000101100; // input=0.75830078125, output=0.860702604419
			11'd777: out = 32'b00000000000000000110111001011101; // input=0.75927734375, output=0.86220192628
			11'd778: out = 32'b00000000000000000110111010001110; // input=0.76025390625, output=0.863703875539
			11'd779: out = 32'b00000000000000000110111010111111; // input=0.76123046875, output=0.865208469465
			11'd780: out = 32'b00000000000000000110111011110001; // input=0.76220703125, output=0.866715725501
			11'd781: out = 32'b00000000000000000110111100100010; // input=0.76318359375, output=0.868225661271
			11'd782: out = 32'b00000000000000000110111101010100; // input=0.76416015625, output=0.869738294579
			11'd783: out = 32'b00000000000000000110111110000101; // input=0.76513671875, output=0.871253643414
			11'd784: out = 32'b00000000000000000110111110110111; // input=0.76611328125, output=0.872771725953
			11'd785: out = 32'b00000000000000000110111111101001; // input=0.76708984375, output=0.874292560562
			11'd786: out = 32'b00000000000000000111000000011011; // input=0.76806640625, output=0.875816165799
			11'd787: out = 32'b00000000000000000111000001001101; // input=0.76904296875, output=0.877342560418
			11'd788: out = 32'b00000000000000000111000001111111; // input=0.77001953125, output=0.878871763373
			11'd789: out = 32'b00000000000000000111000010110001; // input=0.77099609375, output=0.880403793817
			11'd790: out = 32'b00000000000000000111000011100011; // input=0.77197265625, output=0.881938671108
			11'd791: out = 32'b00000000000000000111000100010110; // input=0.77294921875, output=0.883476414811
			11'd792: out = 32'b00000000000000000111000101001000; // input=0.77392578125, output=0.885017044704
			11'd793: out = 32'b00000000000000000111000101111011; // input=0.77490234375, output=0.886560580776
			11'd794: out = 32'b00000000000000000111000110101101; // input=0.77587890625, output=0.888107043235
			11'd795: out = 32'b00000000000000000111000111100000; // input=0.77685546875, output=0.889656452506
			11'd796: out = 32'b00000000000000000111001000010011; // input=0.77783203125, output=0.891208829243
			11'd797: out = 32'b00000000000000000111001001000110; // input=0.77880859375, output=0.892764194322
			11'd798: out = 32'b00000000000000000111001001111001; // input=0.77978515625, output=0.894322568854
			11'd799: out = 32'b00000000000000000111001010101100; // input=0.78076171875, output=0.895883974181
			11'd800: out = 32'b00000000000000000111001011100000; // input=0.78173828125, output=0.897448431885
			11'd801: out = 32'b00000000000000000111001100010011; // input=0.78271484375, output=0.899015963789
			11'd802: out = 32'b00000000000000000111001101000110; // input=0.78369140625, output=0.900586591962
			11'd803: out = 32'b00000000000000000111001101111010; // input=0.78466796875, output=0.902160338722
			11'd804: out = 32'b00000000000000000111001110101110; // input=0.78564453125, output=0.903737226641
			11'd805: out = 32'b00000000000000000111001111100001; // input=0.78662109375, output=0.905317278548
			11'd806: out = 32'b00000000000000000111010000010101; // input=0.78759765625, output=0.906900517533
			11'd807: out = 32'b00000000000000000111010001001001; // input=0.78857421875, output=0.908486966953
			11'd808: out = 32'b00000000000000000111010001111101; // input=0.78955078125, output=0.910076650436
			11'd809: out = 32'b00000000000000000111010010110010; // input=0.79052734375, output=0.911669591883
			11'd810: out = 32'b00000000000000000111010011100110; // input=0.79150390625, output=0.913265815473
			11'd811: out = 32'b00000000000000000111010100011010; // input=0.79248046875, output=0.914865345673
			11'd812: out = 32'b00000000000000000111010101001111; // input=0.79345703125, output=0.916468207233
			11'd813: out = 32'b00000000000000000111010110000011; // input=0.79443359375, output=0.918074425201
			11'd814: out = 32'b00000000000000000111010110111000; // input=0.79541015625, output=0.919684024919
			11'd815: out = 32'b00000000000000000111010111101101; // input=0.79638671875, output=0.921297032036
			11'd816: out = 32'b00000000000000000111011000100010; // input=0.79736328125, output=0.922913472506
			11'd817: out = 32'b00000000000000000111011001010111; // input=0.79833984375, output=0.924533372597
			11'd818: out = 32'b00000000000000000111011010001100; // input=0.79931640625, output=0.926156758898
			11'd819: out = 32'b00000000000000000111011011000010; // input=0.80029296875, output=0.92778365832
			11'd820: out = 32'b00000000000000000111011011110111; // input=0.80126953125, output=0.929414098105
			11'd821: out = 32'b00000000000000000111011100101101; // input=0.80224609375, output=0.931048105828
			11'd822: out = 32'b00000000000000000111011101100010; // input=0.80322265625, output=0.932685709409
			11'd823: out = 32'b00000000000000000111011110011000; // input=0.80419921875, output=0.934326937112
			11'd824: out = 32'b00000000000000000111011111001110; // input=0.80517578125, output=0.935971817557
			11'd825: out = 32'b00000000000000000111100000000100; // input=0.80615234375, output=0.937620379721
			11'd826: out = 32'b00000000000000000111100000111010; // input=0.80712890625, output=0.93927265295
			11'd827: out = 32'b00000000000000000111100001110000; // input=0.80810546875, output=0.940928666959
			11'd828: out = 32'b00000000000000000111100010100111; // input=0.80908203125, output=0.942588451845
			11'd829: out = 32'b00000000000000000111100011011101; // input=0.81005859375, output=0.944252038088
			11'd830: out = 32'b00000000000000000111100100010100; // input=0.81103515625, output=0.945919456565
			11'd831: out = 32'b00000000000000000111100101001011; // input=0.81201171875, output=0.947590738548
			11'd832: out = 32'b00000000000000000111100110000010; // input=0.81298828125, output=0.949265915721
			11'd833: out = 32'b00000000000000000111100110111001; // input=0.81396484375, output=0.95094502018
			11'd834: out = 32'b00000000000000000111100111110000; // input=0.81494140625, output=0.952628084445
			11'd835: out = 32'b00000000000000000111101000100111; // input=0.81591796875, output=0.954315141464
			11'd836: out = 32'b00000000000000000111101001011110; // input=0.81689453125, output=0.956006224626
			11'd837: out = 32'b00000000000000000111101010010110; // input=0.81787109375, output=0.957701367765
			11'd838: out = 32'b00000000000000000111101011001110; // input=0.81884765625, output=0.95940060517
			11'd839: out = 32'b00000000000000000111101100000101; // input=0.81982421875, output=0.961103971595
			11'd840: out = 32'b00000000000000000111101100111101; // input=0.82080078125, output=0.962811502264
			11'd841: out = 32'b00000000000000000111101101110101; // input=0.82177734375, output=0.964523232885
			11'd842: out = 32'b00000000000000000111101110101110; // input=0.82275390625, output=0.966239199654
			11'd843: out = 32'b00000000000000000111101111100110; // input=0.82373046875, output=0.967959439271
			11'd844: out = 32'b00000000000000000111110000011111; // input=0.82470703125, output=0.969683988941
			11'd845: out = 32'b00000000000000000111110001010111; // input=0.82568359375, output=0.971412886393
			11'd846: out = 32'b00000000000000000111110010010000; // input=0.82666015625, output=0.973146169884
			11'd847: out = 32'b00000000000000000111110011001001; // input=0.82763671875, output=0.974883878213
			11'd848: out = 32'b00000000000000000111110100000010; // input=0.82861328125, output=0.976626050731
			11'd849: out = 32'b00000000000000000111110100111011; // input=0.82958984375, output=0.978372727348
			11'd850: out = 32'b00000000000000000111110101110101; // input=0.83056640625, output=0.980123948551
			11'd851: out = 32'b00000000000000000111110110101110; // input=0.83154296875, output=0.981879755413
			11'd852: out = 32'b00000000000000000111110111101000; // input=0.83251953125, output=0.983640189601
			11'd853: out = 32'b00000000000000000111111000100010; // input=0.83349609375, output=0.985405293394
			11'd854: out = 32'b00000000000000000111111001011100; // input=0.83447265625, output=0.987175109694
			11'd855: out = 32'b00000000000000000111111010010110; // input=0.83544921875, output=0.988949682035
			11'd856: out = 32'b00000000000000000111111011010000; // input=0.83642578125, output=0.990729054601
			11'd857: out = 32'b00000000000000000111111100001011; // input=0.83740234375, output=0.992513272239
			11'd858: out = 32'b00000000000000000111111101000101; // input=0.83837890625, output=0.99430238047
			11'd859: out = 32'b00000000000000000111111110000000; // input=0.83935546875, output=0.996096425507
			11'd860: out = 32'b00000000000000000111111110111011; // input=0.84033203125, output=0.997895454266
			11'd861: out = 32'b00000000000000000111111111110110; // input=0.84130859375, output=0.999699514384
			11'd862: out = 32'b00000000000000001000000000110001; // input=0.84228515625, output=1.00150865423
			11'd863: out = 32'b00000000000000001000000001101101; // input=0.84326171875, output=1.00332292294
			11'd864: out = 32'b00000000000000001000000010101001; // input=0.84423828125, output=1.00514237039
			11'd865: out = 32'b00000000000000001000000011100100; // input=0.84521484375, output=1.00696704727
			11'd866: out = 32'b00000000000000001000000100100000; // input=0.84619140625, output=1.00879700506
			11'd867: out = 32'b00000000000000001000000101011100; // input=0.84716796875, output=1.01063229605
			11'd868: out = 32'b00000000000000001000000110011001; // input=0.84814453125, output=1.01247297339
			11'd869: out = 32'b00000000000000001000000111010101; // input=0.84912109375, output=1.01431909107
			11'd870: out = 32'b00000000000000001000001000010010; // input=0.85009765625, output=1.01617070397
			11'd871: out = 32'b00000000000000001000001001001111; // input=0.85107421875, output=1.01802786786
			11'd872: out = 32'b00000000000000001000001010001100; // input=0.85205078125, output=1.01989063942
			11'd873: out = 32'b00000000000000001000001011001001; // input=0.85302734375, output=1.02175907629
			11'd874: out = 32'b00000000000000001000001100000110; // input=0.85400390625, output=1.02363323705
			11'd875: out = 32'b00000000000000001000001101000100; // input=0.85498046875, output=1.02551318129
			11'd876: out = 32'b00000000000000001000001110000010; // input=0.85595703125, output=1.02739896957
			11'd877: out = 32'b00000000000000001000001111000000; // input=0.85693359375, output=1.02929066351
			11'd878: out = 32'b00000000000000001000001111111110; // input=0.85791015625, output=1.03118832579
			11'd879: out = 32'b00000000000000001000010000111100; // input=0.85888671875, output=1.03309202014
			11'd880: out = 32'b00000000000000001000010001111011; // input=0.85986328125, output=1.03500181142
			11'd881: out = 32'b00000000000000001000010010111010; // input=0.86083984375, output=1.03691776563
			11'd882: out = 32'b00000000000000001000010011111001; // input=0.86181640625, output=1.03883994992
			11'd883: out = 32'b00000000000000001000010100111000; // input=0.86279296875, output=1.04076843263
			11'd884: out = 32'b00000000000000001000010101110111; // input=0.86376953125, output=1.04270328333
			11'd885: out = 32'b00000000000000001000010110110111; // input=0.86474609375, output=1.04464457284
			11'd886: out = 32'b00000000000000001000010111110111; // input=0.86572265625, output=1.04659237326
			11'd887: out = 32'b00000000000000001000011000110111; // input=0.86669921875, output=1.04854675801
			11'd888: out = 32'b00000000000000001000011001110111; // input=0.86767578125, output=1.05050780186
			11'd889: out = 32'b00000000000000001000011010111000; // input=0.86865234375, output=1.05247558096
			11'd890: out = 32'b00000000000000001000011011111000; // input=0.86962890625, output=1.0544501729
			11'd891: out = 32'b00000000000000001000011100111001; // input=0.87060546875, output=1.0564316567
			11'd892: out = 32'b00000000000000001000011101111010; // input=0.87158203125, output=1.0584201129
			11'd893: out = 32'b00000000000000001000011110111100; // input=0.87255859375, output=1.06041562356
			11'd894: out = 32'b00000000000000001000011111111101; // input=0.87353515625, output=1.06241827236
			11'd895: out = 32'b00000000000000001000100000111111; // input=0.87451171875, output=1.06442814454
			11'd896: out = 32'b00000000000000001000100010000001; // input=0.87548828125, output=1.06644532706
			11'd897: out = 32'b00000000000000001000100011000100; // input=0.87646484375, output=1.06846990857
			11'd898: out = 32'b00000000000000001000100100000110; // input=0.87744140625, output=1.07050197947
			11'd899: out = 32'b00000000000000001000100101001001; // input=0.87841796875, output=1.07254163199
			11'd900: out = 32'b00000000000000001000100110001100; // input=0.87939453125, output=1.0745889602
			11'd901: out = 32'b00000000000000001000100111001111; // input=0.88037109375, output=1.07664406011
			11'd902: out = 32'b00000000000000001000101000010011; // input=0.88134765625, output=1.07870702967
			11'd903: out = 32'b00000000000000001000101001010111; // input=0.88232421875, output=1.08077796888
			11'd904: out = 32'b00000000000000001000101010011011; // input=0.88330078125, output=1.08285697979
			11'd905: out = 32'b00000000000000001000101011011111; // input=0.88427734375, output=1.08494416663
			11'd906: out = 32'b00000000000000001000101100100100; // input=0.88525390625, output=1.08703963583
			11'd907: out = 32'b00000000000000001000101101101001; // input=0.88623046875, output=1.08914349607
			11'd908: out = 32'b00000000000000001000101110101110; // input=0.88720703125, output=1.09125585841
			11'd909: out = 32'b00000000000000001000101111110100; // input=0.88818359375, output=1.09337683631
			11'd910: out = 32'b00000000000000001000110000111010; // input=0.88916015625, output=1.0955065457
			11'd911: out = 32'b00000000000000001000110010000000; // input=0.89013671875, output=1.0976451051
			11'd912: out = 32'b00000000000000001000110011000110; // input=0.89111328125, output=1.09979263568
			11'd913: out = 32'b00000000000000001000110100001101; // input=0.89208984375, output=1.10194926132
			11'd914: out = 32'b00000000000000001000110101010100; // input=0.89306640625, output=1.10411510871
			11'd915: out = 32'b00000000000000001000110110011011; // input=0.89404296875, output=1.10629030749
			11'd916: out = 32'b00000000000000001000110111100011; // input=0.89501953125, output=1.10847499025
			11'd917: out = 32'b00000000000000001000111000101010; // input=0.89599609375, output=1.1106692927
			11'd918: out = 32'b00000000000000001000111001110011; // input=0.89697265625, output=1.11287335376
			11'd919: out = 32'b00000000000000001000111010111011; // input=0.89794921875, output=1.11508731565
			11'd920: out = 32'b00000000000000001000111100000100; // input=0.89892578125, output=1.117311324
			11'd921: out = 32'b00000000000000001000111101001101; // input=0.89990234375, output=1.11954552799
			11'd922: out = 32'b00000000000000001000111110010111; // input=0.90087890625, output=1.12179008044
			11'd923: out = 32'b00000000000000001000111111100001; // input=0.90185546875, output=1.12404513797
			11'd924: out = 32'b00000000000000001001000000101011; // input=0.90283203125, output=1.1263108611
			11'd925: out = 32'b00000000000000001001000001110110; // input=0.90380859375, output=1.12858741441
			11'd926: out = 32'b00000000000000001001000011000001; // input=0.90478515625, output=1.13087496667
			11'd927: out = 32'b00000000000000001001000100001100; // input=0.90576171875, output=1.13317369102
			11'd928: out = 32'b00000000000000001001000101011000; // input=0.90673828125, output=1.13548376509
			11'd929: out = 32'b00000000000000001001000110100100; // input=0.90771484375, output=1.13780537118
			11'd930: out = 32'b00000000000000001001000111110000; // input=0.90869140625, output=1.14013869645
			11'd931: out = 32'b00000000000000001001001000111101; // input=0.90966796875, output=1.14248393307
			11'd932: out = 32'b00000000000000001001001010001010; // input=0.91064453125, output=1.14484127846
			11'd933: out = 32'b00000000000000001001001011011000; // input=0.91162109375, output=1.14721093543
			11'd934: out = 32'b00000000000000001001001100100110; // input=0.91259765625, output=1.14959311244
			11'd935: out = 32'b00000000000000001001001101110100; // input=0.91357421875, output=1.1519880238
			11'd936: out = 32'b00000000000000001001001111000011; // input=0.91455078125, output=1.1543958899
			11'd937: out = 32'b00000000000000001001010000010011; // input=0.91552734375, output=1.15681693745
			11'd938: out = 32'b00000000000000001001010001100010; // input=0.91650390625, output=1.15925139978
			11'd939: out = 32'b00000000000000001001010010110011; // input=0.91748046875, output=1.16169951703
			11'd940: out = 32'b00000000000000001001010100000011; // input=0.91845703125, output=1.16416153653
			11'd941: out = 32'b00000000000000001001010101010100; // input=0.91943359375, output=1.16663771301
			11'd942: out = 32'b00000000000000001001010110100110; // input=0.92041015625, output=1.16912830899
			11'd943: out = 32'b00000000000000001001010111111000; // input=0.92138671875, output=1.17163359507
			11'd944: out = 32'b00000000000000001001011001001011; // input=0.92236328125, output=1.17415385031
			11'd945: out = 32'b00000000000000001001011010011110; // input=0.92333984375, output=1.17668936258
			11'd946: out = 32'b00000000000000001001011011110001; // input=0.92431640625, output=1.17924042897
			11'd947: out = 32'b00000000000000001001011101000101; // input=0.92529296875, output=1.18180735621
			11'd948: out = 32'b00000000000000001001011110011010; // input=0.92626953125, output=1.1843904611
			11'd949: out = 32'b00000000000000001001011111101111; // input=0.92724609375, output=1.18699007099
			11'd950: out = 32'b00000000000000001001100001000101; // input=0.92822265625, output=1.18960652428
			11'd951: out = 32'b00000000000000001001100010011011; // input=0.92919921875, output=1.19224017094
			11'd952: out = 32'b00000000000000001001100011110010; // input=0.93017578125, output=1.19489137306
			11'd953: out = 32'b00000000000000001001100101001010; // input=0.93115234375, output=1.1975605055
			11'd954: out = 32'b00000000000000001001100110100010; // input=0.93212890625, output=1.20024795643
			11'd955: out = 32'b00000000000000001001100111111010; // input=0.93310546875, output=1.20295412811
			11'd956: out = 32'b00000000000000001001101001010100; // input=0.93408203125, output=1.20567943755
			11'd957: out = 32'b00000000000000001001101010101110; // input=0.93505859375, output=1.20842431728
			11'd958: out = 32'b00000000000000001001101100001000; // input=0.93603515625, output=1.21118921619
			11'd959: out = 32'b00000000000000001001101101100100; // input=0.93701171875, output=1.2139746004
			11'd960: out = 32'b00000000000000001001101110111111; // input=0.93798828125, output=1.21678095422
			11'd961: out = 32'b00000000000000001001110000011100; // input=0.93896484375, output=1.21960878111
			11'd962: out = 32'b00000000000000001001110001111010; // input=0.93994140625, output=1.22245860481
			11'd963: out = 32'b00000000000000001001110011011000; // input=0.94091796875, output=1.22533097047
			11'd964: out = 32'b00000000000000001001110100110111; // input=0.94189453125, output=1.22822644589
			11'd965: out = 32'b00000000000000001001110110010110; // input=0.94287109375, output=1.23114562288
			11'd966: out = 32'b00000000000000001001110111110111; // input=0.94384765625, output=1.23408911871
			11'd967: out = 32'b00000000000000001001111001011000; // input=0.94482421875, output=1.23705757763
			11'd968: out = 32'b00000000000000001001111010111010; // input=0.94580078125, output=1.24005167258
			11'd969: out = 32'b00000000000000001001111100011101; // input=0.94677734375, output=1.24307210702
			11'd970: out = 32'b00000000000000001001111110000001; // input=0.94775390625, output=1.24611961686
			11'd971: out = 32'b00000000000000001001111111100110; // input=0.94873046875, output=1.24919497264
			11'd972: out = 32'b00000000000000001010000001001011; // input=0.94970703125, output=1.25229898181
			11'd973: out = 32'b00000000000000001010000010110010; // input=0.95068359375, output=1.25543249128
			11'd974: out = 32'b00000000000000001010000100011010; // input=0.95166015625, output=1.25859639018
			11'd975: out = 32'b00000000000000001010000110000010; // input=0.95263671875, output=1.26179161284
			11'd976: out = 32'b00000000000000001010000111101100; // input=0.95361328125, output=1.26501914206
			11'd977: out = 32'b00000000000000001010001001010111; // input=0.95458984375, output=1.26828001276
			11'd978: out = 32'b00000000000000001010001011000011; // input=0.95556640625, output=1.27157531586
			11'd979: out = 32'b00000000000000001010001100110000; // input=0.95654296875, output=1.27490620266
			11'd980: out = 32'b00000000000000001010001110011110; // input=0.95751953125, output=1.27827388961
			11'd981: out = 32'b00000000000000001010010000001110; // input=0.95849609375, output=1.28167966359
			11'd982: out = 32'b00000000000000001010010001111111; // input=0.95947265625, output=1.28512488772
			11'd983: out = 32'b00000000000000001010010011110001; // input=0.96044921875, output=1.28861100788
			11'd984: out = 32'b00000000000000001010010101100101; // input=0.96142578125, output=1.2921395599
			11'd985: out = 32'b00000000000000001010010111011010; // input=0.96240234375, output=1.29571217755
			11'd986: out = 32'b00000000000000001010011001010000; // input=0.96337890625, output=1.29933060156
			11'd987: out = 32'b00000000000000001010011011001001; // input=0.96435546875, output=1.30299668967
			11'd988: out = 32'b00000000000000001010011101000010; // input=0.96533203125, output=1.30671242792
			11'd989: out = 32'b00000000000000001010011110111110; // input=0.96630859375, output=1.3104799434
			11'd990: out = 32'b00000000000000001010100000111011; // input=0.96728515625, output=1.31430151869
			11'd991: out = 32'b00000000000000001010100010111010; // input=0.96826171875, output=1.31817960826
			11'd992: out = 32'b00000000000000001010100100111011; // input=0.96923828125, output=1.32211685711
			11'd993: out = 32'b00000000000000001010100110111110; // input=0.97021484375, output=1.32611612215
			11'd994: out = 32'b00000000000000001010101001000011; // input=0.97119140625, output=1.33018049673
			11'd995: out = 32'b00000000000000001010101011001011; // input=0.97216796875, output=1.33431333899
			11'd996: out = 32'b00000000000000001010101101010101; // input=0.97314453125, output=1.33851830468
			11'd997: out = 32'b00000000000000001010101111100001; // input=0.97412109375, output=1.34279938541
			11'd998: out = 32'b00000000000000001010110001110000; // input=0.97509765625, output=1.34716095354
			11'd999: out = 32'b00000000000000001010110100000001; // input=0.97607421875, output=1.35160781497
			11'd1000: out = 32'b00000000000000001010110110010110; // input=0.97705078125, output=1.35614527182
			11'd1001: out = 32'b00000000000000001010111000101110; // input=0.97802734375, output=1.36077919721
			11'd1002: out = 32'b00000000000000001010111011001001; // input=0.97900390625, output=1.36551612523
			11'd1003: out = 32'b00000000000000001010111101101000; // input=0.97998046875, output=1.37036335996
			11'd1004: out = 32'b00000000000000001011000000001011; // input=0.98095703125, output=1.37532910873
			11'd1005: out = 32'b00000000000000001011000010110010; // input=0.98193359375, output=1.38042264672
			11'd1006: out = 32'b00000000000000001011000101011101; // input=0.98291015625, output=1.38565452202
			11'd1007: out = 32'b00000000000000001011001000001101; // input=0.98388671875, output=1.39103681451
			11'd1008: out = 32'b00000000000000001011001011000011; // input=0.98486328125, output=1.39658346647
			11'd1009: out = 32'b00000000000000001011001101111111; // input=0.98583984375, output=1.40231071107
			11'd1010: out = 32'b00000000000000001011010001000001; // input=0.98681640625, output=1.40823763659
			11'd1011: out = 32'b00000000000000001011010100001011; // input=0.98779296875, output=1.41438694293
			11'd1012: out = 32'b00000000000000001011010111011100; // input=0.98876953125, output=1.42078597714
			11'd1013: out = 32'b00000000000000001011011010110111; // input=0.98974609375, output=1.42746818517
			11'd1014: out = 32'b00000000000000001011011110011101; // input=0.99072265625, output=1.43447520447
			11'd1015: out = 32'b00000000000000001011100010001111; // input=0.99169921875, output=1.44185998152
			11'd1016: out = 32'b00000000000000001011100110001111; // input=0.99267578125, output=1.44969160393
			11'd1017: out = 32'b00000000000000001011101010100010; // input=0.99365234375, output=1.45806316311
			11'd1018: out = 32'b00000000000000001011101111001010; // input=0.99462890625, output=1.46710535557
			11'd1019: out = 32'b00000000000000001011110100001111; // input=0.99560546875, output=1.47701196053
			11'd1020: out = 32'b00000000000000001011111001111010; // input=0.99658203125, output=1.48809303047
			11'd1021: out = 32'b00000000000000001100000000011110; // input=0.99755859375, output=1.50090497815
			11'd1022: out = 32'b00000000000000001100001000100010; // input=0.99853515625, output=1.51666312963
			11'd1023: out = 32'b00000000000000001100010100010000; // input=0.99951171875, output=1.53954505509
			11'd1024: out = 32'b10000000000000000000000000010000; // input=-0.00048828125, output=-0.000488281269403
			11'd1025: out = 32'b10000000000000000000000000110000; // input=-0.00146484375, output=-0.00146484427387
			11'd1026: out = 32'b10000000000000000000000001010000; // input=-0.00244140625, output=-0.00244140867533
			11'd1027: out = 32'b10000000000000000000000001110000; // input=-0.00341796875, output=-0.00341797540511
			11'd1028: out = 32'b10000000000000000000000010010000; // input=-0.00439453125, output=-0.00439454539458
			11'd1029: out = 32'b10000000000000000000000010110000; // input=-0.00537109375, output=-0.00537111957513
			11'd1030: out = 32'b10000000000000000000000011010000; // input=-0.00634765625, output=-0.00634769887818
			11'd1031: out = 32'b10000000000000000000000011110000; // input=-0.00732421875, output=-0.0073242842352
			11'd1032: out = 32'b10000000000000000000000100010000; // input=-0.00830078125, output=-0.0083008765777
			11'd1033: out = 32'b10000000000000000000000100110000; // input=-0.00927734375, output=-0.00927747683727
			11'd1034: out = 32'b10000000000000000000000101010000; // input=-0.01025390625, output=-0.0102540859456
			11'd1035: out = 32'b10000000000000000000000101110000; // input=-0.01123046875, output=-0.0112307048343
			11'd1036: out = 32'b10000000000000000000000110010000; // input=-0.01220703125, output=-0.0122073344352
			11'd1037: out = 32'b10000000000000000000000110110000; // input=-0.01318359375, output=-0.0131839756803
			11'd1038: out = 32'b10000000000000000000000111010000; // input=-0.01416015625, output=-0.0141606295016
			11'd1039: out = 32'b10000000000000000000000111110000; // input=-0.01513671875, output=-0.0151372968311
			11'd1040: out = 32'b10000000000000000000001000010000; // input=-0.01611328125, output=-0.016113978601
			11'd1041: out = 32'b10000000000000000000001000110000; // input=-0.01708984375, output=-0.0170906757438
			11'd1042: out = 32'b10000000000000000000001001010000; // input=-0.01806640625, output=-0.0180673891919
			11'd1043: out = 32'b10000000000000000000001001110000; // input=-0.01904296875, output=-0.0190441198779
			11'd1044: out = 32'b10000000000000000000001010010000; // input=-0.02001953125, output=-0.0200208687346
			11'd1045: out = 32'b10000000000000000000001010110000; // input=-0.02099609375, output=-0.0209976366949
			11'd1046: out = 32'b10000000000000000000001011010000; // input=-0.02197265625, output=-0.0219744246919
			11'd1047: out = 32'b10000000000000000000001011110000; // input=-0.02294921875, output=-0.0229512336589
			11'd1048: out = 32'b10000000000000000000001100010000; // input=-0.02392578125, output=-0.0239280645293
			11'd1049: out = 32'b10000000000000000000001100110000; // input=-0.02490234375, output=-0.0249049182366
			11'd1050: out = 32'b10000000000000000000001101010000; // input=-0.02587890625, output=-0.0258817957149
			11'd1051: out = 32'b10000000000000000000001101110000; // input=-0.02685546875, output=-0.026858697898
			11'd1052: out = 32'b10000000000000000000001110010000; // input=-0.02783203125, output=-0.0278356257202
			11'd1053: out = 32'b10000000000000000000001110110000; // input=-0.02880859375, output=-0.028812580116
			11'd1054: out = 32'b10000000000000000000001111010000; // input=-0.02978515625, output=-0.0297895620201
			11'd1055: out = 32'b10000000000000000000001111110000; // input=-0.03076171875, output=-0.0307665723674
			11'd1056: out = 32'b10000000000000000000010000010000; // input=-0.03173828125, output=-0.0317436120931
			11'd1057: out = 32'b10000000000000000000010000110000; // input=-0.03271484375, output=-0.0327206821325
			11'd1058: out = 32'b10000000000000000000010001010000; // input=-0.03369140625, output=-0.0336977834215
			11'd1059: out = 32'b10000000000000000000010001110000; // input=-0.03466796875, output=-0.0346749168959
			11'd1060: out = 32'b10000000000000000000010010010000; // input=-0.03564453125, output=-0.0356520834919
			11'd1061: out = 32'b10000000000000000000010010110000; // input=-0.03662109375, output=-0.0366292841462
			11'd1062: out = 32'b10000000000000000000010011010000; // input=-0.03759765625, output=-0.0376065197954
			11'd1063: out = 32'b10000000000000000000010011110000; // input=-0.03857421875, output=-0.0385837913767
			11'd1064: out = 32'b10000000000000000000010100010000; // input=-0.03955078125, output=-0.0395610998276
			11'd1065: out = 32'b10000000000000000000010100110000; // input=-0.04052734375, output=-0.0405384460857
			11'd1066: out = 32'b10000000000000000000010101010000; // input=-0.04150390625, output=-0.0415158310892
			11'd1067: out = 32'b10000000000000000000010101110000; // input=-0.04248046875, output=-0.0424932557764
			11'd1068: out = 32'b10000000000000000000010110010000; // input=-0.04345703125, output=-0.0434707210861
			11'd1069: out = 32'b10000000000000000000010110110000; // input=-0.04443359375, output=-0.0444482279573
			11'd1070: out = 32'b10000000000000000000010111010001; // input=-0.04541015625, output=-0.0454257773296
			11'd1071: out = 32'b10000000000000000000010111110001; // input=-0.04638671875, output=-0.0464033701426
			11'd1072: out = 32'b10000000000000000000011000010001; // input=-0.04736328125, output=-0.0473810073367
			11'd1073: out = 32'b10000000000000000000011000110001; // input=-0.04833984375, output=-0.0483586898524
			11'd1074: out = 32'b10000000000000000000011001010001; // input=-0.04931640625, output=-0.0493364186307
			11'd1075: out = 32'b10000000000000000000011001110001; // input=-0.05029296875, output=-0.0503141946129
			11'd1076: out = 32'b10000000000000000000011010010001; // input=-0.05126953125, output=-0.0512920187407
			11'd1077: out = 32'b10000000000000000000011010110001; // input=-0.05224609375, output=-0.0522698919565
			11'd1078: out = 32'b10000000000000000000011011010001; // input=-0.05322265625, output=-0.0532478152028
			11'd1079: out = 32'b10000000000000000000011011110001; // input=-0.05419921875, output=-0.0542257894226
			11'd1080: out = 32'b10000000000000000000011100010001; // input=-0.05517578125, output=-0.0552038155595
			11'd1081: out = 32'b10000000000000000000011100110001; // input=-0.05615234375, output=-0.0561818945573
			11'd1082: out = 32'b10000000000000000000011101010001; // input=-0.05712890625, output=-0.0571600273605
			11'd1083: out = 32'b10000000000000000000011101110001; // input=-0.05810546875, output=-0.0581382149139
			11'd1084: out = 32'b10000000000000000000011110010001; // input=-0.05908203125, output=-0.0591164581629
			11'd1085: out = 32'b10000000000000000000011110110001; // input=-0.06005859375, output=-0.0600947580532
			11'd1086: out = 32'b10000000000000000000011111010001; // input=-0.06103515625, output=-0.0610731155313
			11'd1087: out = 32'b10000000000000000000011111110001; // input=-0.06201171875, output=-0.0620515315438
			11'd1088: out = 32'b10000000000000000000100000010001; // input=-0.06298828125, output=-0.0630300070381
			11'd1089: out = 32'b10000000000000000000100000110001; // input=-0.06396484375, output=-0.064008542962
			11'd1090: out = 32'b10000000000000000000100001010001; // input=-0.06494140625, output=-0.064987140264
			11'd1091: out = 32'b10000000000000000000100001110010; // input=-0.06591796875, output=-0.0659657998927
			11'd1092: out = 32'b10000000000000000000100010010010; // input=-0.06689453125, output=-0.0669445227978
			11'd1093: out = 32'b10000000000000000000100010110010; // input=-0.06787109375, output=-0.0679233099292
			11'd1094: out = 32'b10000000000000000000100011010010; // input=-0.06884765625, output=-0.0689021622373
			11'd1095: out = 32'b10000000000000000000100011110010; // input=-0.06982421875, output=-0.0698810806733
			11'd1096: out = 32'b10000000000000000000100100010010; // input=-0.07080078125, output=-0.070860066189
			11'd1097: out = 32'b10000000000000000000100100110010; // input=-0.07177734375, output=-0.0718391197364
			11'd1098: out = 32'b10000000000000000000100101010010; // input=-0.07275390625, output=-0.0728182422686
			11'd1099: out = 32'b10000000000000000000100101110010; // input=-0.07373046875, output=-0.0737974347388
			11'd1100: out = 32'b10000000000000000000100110010010; // input=-0.07470703125, output=-0.0747766981013
			11'd1101: out = 32'b10000000000000000000100110110010; // input=-0.07568359375, output=-0.0757560333106
			11'd1102: out = 32'b10000000000000000000100111010010; // input=-0.07666015625, output=-0.0767354413221
			11'd1103: out = 32'b10000000000000000000100111110011; // input=-0.07763671875, output=-0.0777149230917
			11'd1104: out = 32'b10000000000000000000101000010011; // input=-0.07861328125, output=-0.0786944795761
			11'd1105: out = 32'b10000000000000000000101000110011; // input=-0.07958984375, output=-0.0796741117323
			11'd1106: out = 32'b10000000000000000000101001010011; // input=-0.08056640625, output=-0.0806538205183
			11'd1107: out = 32'b10000000000000000000101001110011; // input=-0.08154296875, output=-0.0816336068927
			11'd1108: out = 32'b10000000000000000000101010010011; // input=-0.08251953125, output=-0.0826134718148
			11'd1109: out = 32'b10000000000000000000101010110011; // input=-0.08349609375, output=-0.0835934162443
			11'd1110: out = 32'b10000000000000000000101011010011; // input=-0.08447265625, output=-0.084573441142
			11'd1111: out = 32'b10000000000000000000101011110011; // input=-0.08544921875, output=-0.0855535474692
			11'd1112: out = 32'b10000000000000000000101100010100; // input=-0.08642578125, output=-0.086533736188
			11'd1113: out = 32'b10000000000000000000101100110100; // input=-0.08740234375, output=-0.087514008261
			11'd1114: out = 32'b10000000000000000000101101010100; // input=-0.08837890625, output=-0.0884943646517
			11'd1115: out = 32'b10000000000000000000101101110100; // input=-0.08935546875, output=-0.0894748063244
			11'd1116: out = 32'b10000000000000000000101110010100; // input=-0.09033203125, output=-0.0904553342441
			11'd1117: out = 32'b10000000000000000000101110110100; // input=-0.09130859375, output=-0.0914359493765
			11'd1118: out = 32'b10000000000000000000101111010100; // input=-0.09228515625, output=-0.0924166526881
			11'd1119: out = 32'b10000000000000000000101111110100; // input=-0.09326171875, output=-0.0933974451461
			11'd1120: out = 32'b10000000000000000000110000010101; // input=-0.09423828125, output=-0.0943783277186
			11'd1121: out = 32'b10000000000000000000110000110101; // input=-0.09521484375, output=-0.0953593013745
			11'd1122: out = 32'b10000000000000000000110001010101; // input=-0.09619140625, output=-0.0963403670833
			11'd1123: out = 32'b10000000000000000000110001110101; // input=-0.09716796875, output=-0.0973215258156
			11'd1124: out = 32'b10000000000000000000110010010101; // input=-0.09814453125, output=-0.0983027785426
			11'd1125: out = 32'b10000000000000000000110010110101; // input=-0.09912109375, output=-0.0992841262364
			11'd1126: out = 32'b10000000000000000000110011010110; // input=-0.10009765625, output=-0.10026556987
			11'd1127: out = 32'b10000000000000000000110011110110; // input=-0.10107421875, output=-0.101247110417
			11'd1128: out = 32'b10000000000000000000110100010110; // input=-0.10205078125, output=-0.102228748852
			11'd1129: out = 32'b10000000000000000000110100110110; // input=-0.10302734375, output=-0.103210486151
			11'd1130: out = 32'b10000000000000000000110101010110; // input=-0.10400390625, output=-0.10419232329
			11'd1131: out = 32'b10000000000000000000110101110110; // input=-0.10498046875, output=-0.105174261246
			11'd1132: out = 32'b10000000000000000000110110010111; // input=-0.10595703125, output=-0.106156300998
			11'd1133: out = 32'b10000000000000000000110110110111; // input=-0.10693359375, output=-0.107138443524
			11'd1134: out = 32'b10000000000000000000110111010111; // input=-0.10791015625, output=-0.108120689804
			11'd1135: out = 32'b10000000000000000000110111110111; // input=-0.10888671875, output=-0.10910304082
			11'd1136: out = 32'b10000000000000000000111000010111; // input=-0.10986328125, output=-0.110085497553
			11'd1137: out = 32'b10000000000000000000111000110111; // input=-0.11083984375, output=-0.111068060986
			11'd1138: out = 32'b10000000000000000000111001011000; // input=-0.11181640625, output=-0.112050732102
			11'd1139: out = 32'b10000000000000000000111001111000; // input=-0.11279296875, output=-0.113033511886
			11'd1140: out = 32'b10000000000000000000111010011000; // input=-0.11376953125, output=-0.114016401324
			11'd1141: out = 32'b10000000000000000000111010111000; // input=-0.11474609375, output=-0.114999401402
			11'd1142: out = 32'b10000000000000000000111011011001; // input=-0.11572265625, output=-0.115982513109
			11'd1143: out = 32'b10000000000000000000111011111001; // input=-0.11669921875, output=-0.116965737431
			11'd1144: out = 32'b10000000000000000000111100011001; // input=-0.11767578125, output=-0.11794907536
			11'd1145: out = 32'b10000000000000000000111100111001; // input=-0.11865234375, output=-0.118932527885
			11'd1146: out = 32'b10000000000000000000111101011001; // input=-0.11962890625, output=-0.119916095998
			11'd1147: out = 32'b10000000000000000000111101111010; // input=-0.12060546875, output=-0.120899780692
			11'd1148: out = 32'b10000000000000000000111110011010; // input=-0.12158203125, output=-0.12188358296
			11'd1149: out = 32'b10000000000000000000111110111010; // input=-0.12255859375, output=-0.122867503798
			11'd1150: out = 32'b10000000000000000000111111011010; // input=-0.12353515625, output=-0.1238515442
			11'd1151: out = 32'b10000000000000000000111111111011; // input=-0.12451171875, output=-0.124835705164
			11'd1152: out = 32'b10000000000000000001000000011011; // input=-0.12548828125, output=-0.125819987687
			11'd1153: out = 32'b10000000000000000001000000111011; // input=-0.12646484375, output=-0.126804392769
			11'd1154: out = 32'b10000000000000000001000001011011; // input=-0.12744140625, output=-0.12778892141
			11'd1155: out = 32'b10000000000000000001000001111100; // input=-0.12841796875, output=-0.12877357461
			11'd1156: out = 32'b10000000000000000001000010011100; // input=-0.12939453125, output=-0.129758353373
			11'd1157: out = 32'b10000000000000000001000010111100; // input=-0.13037109375, output=-0.130743258701
			11'd1158: out = 32'b10000000000000000001000011011100; // input=-0.13134765625, output=-0.1317282916
			11'd1159: out = 32'b10000000000000000001000011111101; // input=-0.13232421875, output=-0.132713453074
			11'd1160: out = 32'b10000000000000000001000100011101; // input=-0.13330078125, output=-0.133698744131
			11'd1161: out = 32'b10000000000000000001000100111101; // input=-0.13427734375, output=-0.134684165779
			11'd1162: out = 32'b10000000000000000001000101011110; // input=-0.13525390625, output=-0.135669719027
			11'd1163: out = 32'b10000000000000000001000101111110; // input=-0.13623046875, output=-0.136655404886
			11'd1164: out = 32'b10000000000000000001000110011110; // input=-0.13720703125, output=-0.137641224367
			11'd1165: out = 32'b10000000000000000001000110111111; // input=-0.13818359375, output=-0.138627178482
			11'd1166: out = 32'b10000000000000000001000111011111; // input=-0.13916015625, output=-0.139613268246
			11'd1167: out = 32'b10000000000000000001000111111111; // input=-0.14013671875, output=-0.140599494675
			11'd1168: out = 32'b10000000000000000001001000011111; // input=-0.14111328125, output=-0.141585858784
			11'd1169: out = 32'b10000000000000000001001001000000; // input=-0.14208984375, output=-0.142572361592
			11'd1170: out = 32'b10000000000000000001001001100000; // input=-0.14306640625, output=-0.143559004117
			11'd1171: out = 32'b10000000000000000001001010000000; // input=-0.14404296875, output=-0.144545787379
			11'd1172: out = 32'b10000000000000000001001010100001; // input=-0.14501953125, output=-0.145532712401
			11'd1173: out = 32'b10000000000000000001001011000001; // input=-0.14599609375, output=-0.146519780204
			11'd1174: out = 32'b10000000000000000001001011100010; // input=-0.14697265625, output=-0.147506991814
			11'd1175: out = 32'b10000000000000000001001100000010; // input=-0.14794921875, output=-0.148494348255
			11'd1176: out = 32'b10000000000000000001001100100010; // input=-0.14892578125, output=-0.149481850554
			11'd1177: out = 32'b10000000000000000001001101000011; // input=-0.14990234375, output=-0.15046949974
			11'd1178: out = 32'b10000000000000000001001101100011; // input=-0.15087890625, output=-0.151457296841
			11'd1179: out = 32'b10000000000000000001001110000011; // input=-0.15185546875, output=-0.152445242889
			11'd1180: out = 32'b10000000000000000001001110100100; // input=-0.15283203125, output=-0.153433338915
			11'd1181: out = 32'b10000000000000000001001111000100; // input=-0.15380859375, output=-0.154421585953
			11'd1182: out = 32'b10000000000000000001001111100100; // input=-0.15478515625, output=-0.155409985038
			11'd1183: out = 32'b10000000000000000001010000000101; // input=-0.15576171875, output=-0.156398537206
			11'd1184: out = 32'b10000000000000000001010000100101; // input=-0.15673828125, output=-0.157387243495
			11'd1185: out = 32'b10000000000000000001010001000110; // input=-0.15771484375, output=-0.158376104944
			11'd1186: out = 32'b10000000000000000001010001100110; // input=-0.15869140625, output=-0.159365122593
			11'd1187: out = 32'b10000000000000000001010010000110; // input=-0.15966796875, output=-0.160354297484
			11'd1188: out = 32'b10000000000000000001010010100111; // input=-0.16064453125, output=-0.161343630661
			11'd1189: out = 32'b10000000000000000001010011000111; // input=-0.16162109375, output=-0.162333123168
			11'd1190: out = 32'b10000000000000000001010011101000; // input=-0.16259765625, output=-0.163322776052
			11'd1191: out = 32'b10000000000000000001010100001000; // input=-0.16357421875, output=-0.16431259036
			11'd1192: out = 32'b10000000000000000001010100101001; // input=-0.16455078125, output=-0.165302567142
			11'd1193: out = 32'b10000000000000000001010101001001; // input=-0.16552734375, output=-0.166292707448
			11'd1194: out = 32'b10000000000000000001010101101010; // input=-0.16650390625, output=-0.167283012331
			11'd1195: out = 32'b10000000000000000001010110001010; // input=-0.16748046875, output=-0.168273482845
			11'd1196: out = 32'b10000000000000000001010110101010; // input=-0.16845703125, output=-0.169264120044
			11'd1197: out = 32'b10000000000000000001010111001011; // input=-0.16943359375, output=-0.170254924986
			11'd1198: out = 32'b10000000000000000001010111101011; // input=-0.17041015625, output=-0.171245898729
			11'd1199: out = 32'b10000000000000000001011000001100; // input=-0.17138671875, output=-0.172237042333
			11'd1200: out = 32'b10000000000000000001011000101100; // input=-0.17236328125, output=-0.173228356859
			11'd1201: out = 32'b10000000000000000001011001001101; // input=-0.17333984375, output=-0.174219843372
			11'd1202: out = 32'b10000000000000000001011001101101; // input=-0.17431640625, output=-0.175211502934
			11'd1203: out = 32'b10000000000000000001011010001110; // input=-0.17529296875, output=-0.176203336613
			11'd1204: out = 32'b10000000000000000001011010101110; // input=-0.17626953125, output=-0.177195345477
			11'd1205: out = 32'b10000000000000000001011011001111; // input=-0.17724609375, output=-0.178187530595
			11'd1206: out = 32'b10000000000000000001011011101111; // input=-0.17822265625, output=-0.179179893039
			11'd1207: out = 32'b10000000000000000001011100010000; // input=-0.17919921875, output=-0.180172433881
			11'd1208: out = 32'b10000000000000000001011100110000; // input=-0.18017578125, output=-0.181165154197
			11'd1209: out = 32'b10000000000000000001011101010001; // input=-0.18115234375, output=-0.182158055061
			11'd1210: out = 32'b10000000000000000001011101110001; // input=-0.18212890625, output=-0.183151137553
			11'd1211: out = 32'b10000000000000000001011110010010; // input=-0.18310546875, output=-0.184144402751
			11'd1212: out = 32'b10000000000000000001011110110011; // input=-0.18408203125, output=-0.185137851738
			11'd1213: out = 32'b10000000000000000001011111010011; // input=-0.18505859375, output=-0.186131485596
			11'd1214: out = 32'b10000000000000000001011111110100; // input=-0.18603515625, output=-0.187125305409
			11'd1215: out = 32'b10000000000000000001100000010100; // input=-0.18701171875, output=-0.188119312266
			11'd1216: out = 32'b10000000000000000001100000110101; // input=-0.18798828125, output=-0.189113507254
			11'd1217: out = 32'b10000000000000000001100001010101; // input=-0.18896484375, output=-0.190107891462
			11'd1218: out = 32'b10000000000000000001100001110110; // input=-0.18994140625, output=-0.191102465984
			11'd1219: out = 32'b10000000000000000001100010010111; // input=-0.19091796875, output=-0.192097231912
			11'd1220: out = 32'b10000000000000000001100010110111; // input=-0.19189453125, output=-0.193092190343
			11'd1221: out = 32'b10000000000000000001100011011000; // input=-0.19287109375, output=-0.194087342373
			11'd1222: out = 32'b10000000000000000001100011111000; // input=-0.19384765625, output=-0.195082689101
			11'd1223: out = 32'b10000000000000000001100100011001; // input=-0.19482421875, output=-0.19607823163
			11'd1224: out = 32'b10000000000000000001100100111010; // input=-0.19580078125, output=-0.19707397106
			11'd1225: out = 32'b10000000000000000001100101011010; // input=-0.19677734375, output=-0.198069908498
			11'd1226: out = 32'b10000000000000000001100101111011; // input=-0.19775390625, output=-0.19906604505
			11'd1227: out = 32'b10000000000000000001100110011100; // input=-0.19873046875, output=-0.200062381825
			11'd1228: out = 32'b10000000000000000001100110111100; // input=-0.19970703125, output=-0.201058919932
			11'd1229: out = 32'b10000000000000000001100111011101; // input=-0.20068359375, output=-0.202055660484
			11'd1230: out = 32'b10000000000000000001100111111110; // input=-0.20166015625, output=-0.203052604596
			11'd1231: out = 32'b10000000000000000001101000011110; // input=-0.20263671875, output=-0.204049753384
			11'd1232: out = 32'b10000000000000000001101000111111; // input=-0.20361328125, output=-0.205047107966
			11'd1233: out = 32'b10000000000000000001101001100000; // input=-0.20458984375, output=-0.206044669461
			11'd1234: out = 32'b10000000000000000001101010000000; // input=-0.20556640625, output=-0.207042438993
			11'd1235: out = 32'b10000000000000000001101010100001; // input=-0.20654296875, output=-0.208040417685
			11'd1236: out = 32'b10000000000000000001101011000010; // input=-0.20751953125, output=-0.209038606664
			11'd1237: out = 32'b10000000000000000001101011100010; // input=-0.20849609375, output=-0.210037007058
			11'd1238: out = 32'b10000000000000000001101100000011; // input=-0.20947265625, output=-0.211035619996
			11'd1239: out = 32'b10000000000000000001101100100100; // input=-0.21044921875, output=-0.212034446612
			11'd1240: out = 32'b10000000000000000001101101000101; // input=-0.21142578125, output=-0.21303348804
			11'd1241: out = 32'b10000000000000000001101101100101; // input=-0.21240234375, output=-0.214032745416
			11'd1242: out = 32'b10000000000000000001101110000110; // input=-0.21337890625, output=-0.215032219878
			11'd1243: out = 32'b10000000000000000001101110100111; // input=-0.21435546875, output=-0.216031912567
			11'd1244: out = 32'b10000000000000000001101111001000; // input=-0.21533203125, output=-0.217031824626
			11'd1245: out = 32'b10000000000000000001101111101000; // input=-0.21630859375, output=-0.218031957201
			11'd1246: out = 32'b10000000000000000001110000001001; // input=-0.21728515625, output=-0.219032311437
			11'd1247: out = 32'b10000000000000000001110000101010; // input=-0.21826171875, output=-0.220032888484
			11'd1248: out = 32'b10000000000000000001110001001011; // input=-0.21923828125, output=-0.221033689493
			11'd1249: out = 32'b10000000000000000001110001101100; // input=-0.22021484375, output=-0.222034715618
			11'd1250: out = 32'b10000000000000000001110010001100; // input=-0.22119140625, output=-0.223035968015
			11'd1251: out = 32'b10000000000000000001110010101101; // input=-0.22216796875, output=-0.224037447841
			11'd1252: out = 32'b10000000000000000001110011001110; // input=-0.22314453125, output=-0.225039156258
			11'd1253: out = 32'b10000000000000000001110011101111; // input=-0.22412109375, output=-0.226041094426
			11'd1254: out = 32'b10000000000000000001110100010000; // input=-0.22509765625, output=-0.227043263512
			11'd1255: out = 32'b10000000000000000001110100110001; // input=-0.22607421875, output=-0.228045664681
			11'd1256: out = 32'b10000000000000000001110101010001; // input=-0.22705078125, output=-0.229048299103
			11'd1257: out = 32'b10000000000000000001110101110010; // input=-0.22802734375, output=-0.23005116795
			11'd1258: out = 32'b10000000000000000001110110010011; // input=-0.22900390625, output=-0.231054272395
			11'd1259: out = 32'b10000000000000000001110110110100; // input=-0.22998046875, output=-0.232057613615
			11'd1260: out = 32'b10000000000000000001110111010101; // input=-0.23095703125, output=-0.233061192788
			11'd1261: out = 32'b10000000000000000001110111110110; // input=-0.23193359375, output=-0.234065011095
			11'd1262: out = 32'b10000000000000000001111000010111; // input=-0.23291015625, output=-0.23506906972
			11'd1263: out = 32'b10000000000000000001111000111000; // input=-0.23388671875, output=-0.236073369847
			11'd1264: out = 32'b10000000000000000001111001011001; // input=-0.23486328125, output=-0.237077912665
			11'd1265: out = 32'b10000000000000000001111001111001; // input=-0.23583984375, output=-0.238082699365
			11'd1266: out = 32'b10000000000000000001111010011010; // input=-0.23681640625, output=-0.239087731139
			11'd1267: out = 32'b10000000000000000001111010111011; // input=-0.23779296875, output=-0.240093009183
			11'd1268: out = 32'b10000000000000000001111011011100; // input=-0.23876953125, output=-0.241098534694
			11'd1269: out = 32'b10000000000000000001111011111101; // input=-0.23974609375, output=-0.242104308872
			11'd1270: out = 32'b10000000000000000001111100011110; // input=-0.24072265625, output=-0.243110332922
			11'd1271: out = 32'b10000000000000000001111100111111; // input=-0.24169921875, output=-0.244116608046
			11'd1272: out = 32'b10000000000000000001111101100000; // input=-0.24267578125, output=-0.245123135455
			11'd1273: out = 32'b10000000000000000001111110000001; // input=-0.24365234375, output=-0.246129916357
			11'd1274: out = 32'b10000000000000000001111110100010; // input=-0.24462890625, output=-0.247136951966
			11'd1275: out = 32'b10000000000000000001111111000011; // input=-0.24560546875, output=-0.248144243497
			11'd1276: out = 32'b10000000000000000001111111100100; // input=-0.24658203125, output=-0.249151792168
			11'd1277: out = 32'b10000000000000000010000000000101; // input=-0.24755859375, output=-0.2501595992
			11'd1278: out = 32'b10000000000000000010000000100110; // input=-0.24853515625, output=-0.251167665816
			11'd1279: out = 32'b10000000000000000010000001000111; // input=-0.24951171875, output=-0.252175993242
			11'd1280: out = 32'b10000000000000000010000001101000; // input=-0.25048828125, output=-0.253184582706
			11'd1281: out = 32'b10000000000000000010000010001001; // input=-0.25146484375, output=-0.25419343544
			11'd1282: out = 32'b10000000000000000010000010101010; // input=-0.25244140625, output=-0.255202552678
			11'd1283: out = 32'b10000000000000000010000011001100; // input=-0.25341796875, output=-0.256211935655
			11'd1284: out = 32'b10000000000000000010000011101101; // input=-0.25439453125, output=-0.257221585612
			11'd1285: out = 32'b10000000000000000010000100001110; // input=-0.25537109375, output=-0.25823150379
			11'd1286: out = 32'b10000000000000000010000100101111; // input=-0.25634765625, output=-0.259241691435
			11'd1287: out = 32'b10000000000000000010000101010000; // input=-0.25732421875, output=-0.260252149793
			11'd1288: out = 32'b10000000000000000010000101110001; // input=-0.25830078125, output=-0.261262880115
			11'd1289: out = 32'b10000000000000000010000110010010; // input=-0.25927734375, output=-0.262273883654
			11'd1290: out = 32'b10000000000000000010000110110011; // input=-0.26025390625, output=-0.263285161666
			11'd1291: out = 32'b10000000000000000010000111010100; // input=-0.26123046875, output=-0.26429671541
			11'd1292: out = 32'b10000000000000000010000111110110; // input=-0.26220703125, output=-0.265308546147
			11'd1293: out = 32'b10000000000000000010001000010111; // input=-0.26318359375, output=-0.266320655141
			11'd1294: out = 32'b10000000000000000010001000111000; // input=-0.26416015625, output=-0.267333043661
			11'd1295: out = 32'b10000000000000000010001001011001; // input=-0.26513671875, output=-0.268345712975
			11'd1296: out = 32'b10000000000000000010001001111010; // input=-0.26611328125, output=-0.269358664358
			11'd1297: out = 32'b10000000000000000010001010011100; // input=-0.26708984375, output=-0.270371899086
			11'd1298: out = 32'b10000000000000000010001010111101; // input=-0.26806640625, output=-0.271385418436
			11'd1299: out = 32'b10000000000000000010001011011110; // input=-0.26904296875, output=-0.272399223693
			11'd1300: out = 32'b10000000000000000010001011111111; // input=-0.27001953125, output=-0.273413316139
			11'd1301: out = 32'b10000000000000000010001100100000; // input=-0.27099609375, output=-0.274427697064
			11'd1302: out = 32'b10000000000000000010001101000010; // input=-0.27197265625, output=-0.275442367758
			11'd1303: out = 32'b10000000000000000010001101100011; // input=-0.27294921875, output=-0.276457329516
			11'd1304: out = 32'b10000000000000000010001110000100; // input=-0.27392578125, output=-0.277472583634
			11'd1305: out = 32'b10000000000000000010001110100101; // input=-0.27490234375, output=-0.278488131412
			11'd1306: out = 32'b10000000000000000010001111000111; // input=-0.27587890625, output=-0.279503974155
			11'd1307: out = 32'b10000000000000000010001111101000; // input=-0.27685546875, output=-0.280520113167
			11'd1308: out = 32'b10000000000000000010010000001001; // input=-0.27783203125, output=-0.28153654976
			11'd1309: out = 32'b10000000000000000010010000101011; // input=-0.27880859375, output=-0.282553285244
			11'd1310: out = 32'b10000000000000000010010001001100; // input=-0.27978515625, output=-0.283570320937
			11'd1311: out = 32'b10000000000000000010010001101101; // input=-0.28076171875, output=-0.284587658157
			11'd1312: out = 32'b10000000000000000010010010001111; // input=-0.28173828125, output=-0.285605298226
			11'd1313: out = 32'b10000000000000000010010010110000; // input=-0.28271484375, output=-0.28662324247
			11'd1314: out = 32'b10000000000000000010010011010001; // input=-0.28369140625, output=-0.287641492218
			11'd1315: out = 32'b10000000000000000010010011110011; // input=-0.28466796875, output=-0.288660048801
			11'd1316: out = 32'b10000000000000000010010100010100; // input=-0.28564453125, output=-0.289678913555
			11'd1317: out = 32'b10000000000000000010010100110110; // input=-0.28662109375, output=-0.290698087817
			11'd1318: out = 32'b10000000000000000010010101010111; // input=-0.28759765625, output=-0.291717572931
			11'd1319: out = 32'b10000000000000000010010101111000; // input=-0.28857421875, output=-0.292737370241
			11'd1320: out = 32'b10000000000000000010010110011010; // input=-0.28955078125, output=-0.293757481095
			11'd1321: out = 32'b10000000000000000010010110111011; // input=-0.29052734375, output=-0.294777906847
			11'd1322: out = 32'b10000000000000000010010111011101; // input=-0.29150390625, output=-0.29579864885
			11'd1323: out = 32'b10000000000000000010010111111110; // input=-0.29248046875, output=-0.296819708463
			11'd1324: out = 32'b10000000000000000010011000100000; // input=-0.29345703125, output=-0.29784108705
			11'd1325: out = 32'b10000000000000000010011001000001; // input=-0.29443359375, output=-0.298862785975
			11'd1326: out = 32'b10000000000000000010011001100011; // input=-0.29541015625, output=-0.299884806608
			11'd1327: out = 32'b10000000000000000010011010000100; // input=-0.29638671875, output=-0.300907150321
			11'd1328: out = 32'b10000000000000000010011010100110; // input=-0.29736328125, output=-0.30192981849
			11'd1329: out = 32'b10000000000000000010011011000111; // input=-0.29833984375, output=-0.302952812495
			11'd1330: out = 32'b10000000000000000010011011101001; // input=-0.29931640625, output=-0.30397613372
			11'd1331: out = 32'b10000000000000000010011100001010; // input=-0.30029296875, output=-0.304999783551
			11'd1332: out = 32'b10000000000000000010011100101100; // input=-0.30126953125, output=-0.306023763378
			11'd1333: out = 32'b10000000000000000010011101001101; // input=-0.30224609375, output=-0.307048074597
			11'd1334: out = 32'b10000000000000000010011101101111; // input=-0.30322265625, output=-0.308072718603
			11'd1335: out = 32'b10000000000000000010011110010001; // input=-0.30419921875, output=-0.309097696799
			11'd1336: out = 32'b10000000000000000010011110110010; // input=-0.30517578125, output=-0.310123010591
			11'd1337: out = 32'b10000000000000000010011111010100; // input=-0.30615234375, output=-0.311148661385
			11'd1338: out = 32'b10000000000000000010011111110101; // input=-0.30712890625, output=-0.312174650596
			11'd1339: out = 32'b10000000000000000010100000010111; // input=-0.30810546875, output=-0.31320097964
			11'd1340: out = 32'b10000000000000000010100000111001; // input=-0.30908203125, output=-0.314227649936
			11'd1341: out = 32'b10000000000000000010100001011010; // input=-0.31005859375, output=-0.315254662909
			11'd1342: out = 32'b10000000000000000010100001111100; // input=-0.31103515625, output=-0.316282019985
			11'd1343: out = 32'b10000000000000000010100010011110; // input=-0.31201171875, output=-0.317309722597
			11'd1344: out = 32'b10000000000000000010100010111111; // input=-0.31298828125, output=-0.318337772181
			11'd1345: out = 32'b10000000000000000010100011100001; // input=-0.31396484375, output=-0.319366170175
			11'd1346: out = 32'b10000000000000000010100100000011; // input=-0.31494140625, output=-0.320394918022
			11'd1347: out = 32'b10000000000000000010100100100100; // input=-0.31591796875, output=-0.32142401717
			11'd1348: out = 32'b10000000000000000010100101000110; // input=-0.31689453125, output=-0.32245346907
			11'd1349: out = 32'b10000000000000000010100101101000; // input=-0.31787109375, output=-0.323483275177
			11'd1350: out = 32'b10000000000000000010100110001010; // input=-0.31884765625, output=-0.32451343695
			11'd1351: out = 32'b10000000000000000010100110101011; // input=-0.31982421875, output=-0.325543955852
			11'd1352: out = 32'b10000000000000000010100111001101; // input=-0.32080078125, output=-0.326574833351
			11'd1353: out = 32'b10000000000000000010100111101111; // input=-0.32177734375, output=-0.327606070917
			11'd1354: out = 32'b10000000000000000010101000010001; // input=-0.32275390625, output=-0.328637670026
			11'd1355: out = 32'b10000000000000000010101000110011; // input=-0.32373046875, output=-0.329669632158
			11'd1356: out = 32'b10000000000000000010101001010100; // input=-0.32470703125, output=-0.330701958797
			11'd1357: out = 32'b10000000000000000010101001110110; // input=-0.32568359375, output=-0.331734651429
			11'd1358: out = 32'b10000000000000000010101010011000; // input=-0.32666015625, output=-0.332767711548
			11'd1359: out = 32'b10000000000000000010101010111010; // input=-0.32763671875, output=-0.333801140649
			11'd1360: out = 32'b10000000000000000010101011011100; // input=-0.32861328125, output=-0.334834940233
			11'd1361: out = 32'b10000000000000000010101011111110; // input=-0.32958984375, output=-0.335869111804
			11'd1362: out = 32'b10000000000000000010101100100000; // input=-0.33056640625, output=-0.336903656873
			11'd1363: out = 32'b10000000000000000010101101000010; // input=-0.33154296875, output=-0.337938576951
			11'd1364: out = 32'b10000000000000000010101101100011; // input=-0.33251953125, output=-0.338973873558
			11'd1365: out = 32'b10000000000000000010101110000101; // input=-0.33349609375, output=-0.340009548215
			11'd1366: out = 32'b10000000000000000010101110100111; // input=-0.33447265625, output=-0.341045602449
			11'd1367: out = 32'b10000000000000000010101111001001; // input=-0.33544921875, output=-0.34208203779
			11'd1368: out = 32'b10000000000000000010101111101011; // input=-0.33642578125, output=-0.343118855775
			11'd1369: out = 32'b10000000000000000010110000001101; // input=-0.33740234375, output=-0.344156057942
			11'd1370: out = 32'b10000000000000000010110000101111; // input=-0.33837890625, output=-0.345193645838
			11'd1371: out = 32'b10000000000000000010110001010001; // input=-0.33935546875, output=-0.346231621009
			11'd1372: out = 32'b10000000000000000010110001110011; // input=-0.34033203125, output=-0.347269985011
			11'd1373: out = 32'b10000000000000000010110010010101; // input=-0.34130859375, output=-0.348308739401
			11'd1374: out = 32'b10000000000000000010110010110111; // input=-0.34228515625, output=-0.349347885742
			11'd1375: out = 32'b10000000000000000010110011011001; // input=-0.34326171875, output=-0.350387425601
			11'd1376: out = 32'b10000000000000000010110011111100; // input=-0.34423828125, output=-0.351427360551
			11'd1377: out = 32'b10000000000000000010110100011110; // input=-0.34521484375, output=-0.352467692167
			11'd1378: out = 32'b10000000000000000010110101000000; // input=-0.34619140625, output=-0.353508422032
			11'd1379: out = 32'b10000000000000000010110101100010; // input=-0.34716796875, output=-0.354549551733
			11'd1380: out = 32'b10000000000000000010110110000100; // input=-0.34814453125, output=-0.355591082858
			11'd1381: out = 32'b10000000000000000010110110100110; // input=-0.34912109375, output=-0.356633017006
			11'd1382: out = 32'b10000000000000000010110111001000; // input=-0.35009765625, output=-0.357675355776
			11'd1383: out = 32'b10000000000000000010110111101010; // input=-0.35107421875, output=-0.358718100774
			11'd1384: out = 32'b10000000000000000010111000001101; // input=-0.35205078125, output=-0.359761253611
			11'd1385: out = 32'b10000000000000000010111000101111; // input=-0.35302734375, output=-0.360804815901
			11'd1386: out = 32'b10000000000000000010111001010001; // input=-0.35400390625, output=-0.361848789265
			11'd1387: out = 32'b10000000000000000010111001110011; // input=-0.35498046875, output=-0.362893175329
			11'd1388: out = 32'b10000000000000000010111010010110; // input=-0.35595703125, output=-0.363937975722
			11'd1389: out = 32'b10000000000000000010111010111000; // input=-0.35693359375, output=-0.364983192081
			11'd1390: out = 32'b10000000000000000010111011011010; // input=-0.35791015625, output=-0.366028826045
			11'd1391: out = 32'b10000000000000000010111011111100; // input=-0.35888671875, output=-0.367074879261
			11'd1392: out = 32'b10000000000000000010111100011111; // input=-0.35986328125, output=-0.368121353378
			11'd1393: out = 32'b10000000000000000010111101000001; // input=-0.36083984375, output=-0.369168250053
			11'd1394: out = 32'b10000000000000000010111101100011; // input=-0.36181640625, output=-0.370215570947
			11'd1395: out = 32'b10000000000000000010111110000110; // input=-0.36279296875, output=-0.371263317726
			11'd1396: out = 32'b10000000000000000010111110101000; // input=-0.36376953125, output=-0.372311492062
			11'd1397: out = 32'b10000000000000000010111111001010; // input=-0.36474609375, output=-0.373360095631
			11'd1398: out = 32'b10000000000000000010111111101101; // input=-0.36572265625, output=-0.374409130116
			11'd1399: out = 32'b10000000000000000011000000001111; // input=-0.36669921875, output=-0.375458597205
			11'd1400: out = 32'b10000000000000000011000000110001; // input=-0.36767578125, output=-0.37650849859
			11'd1401: out = 32'b10000000000000000011000001010100; // input=-0.36865234375, output=-0.377558835969
			11'd1402: out = 32'b10000000000000000011000001110110; // input=-0.36962890625, output=-0.378609611047
			11'd1403: out = 32'b10000000000000000011000010011001; // input=-0.37060546875, output=-0.379660825532
			11'd1404: out = 32'b10000000000000000011000010111011; // input=-0.37158203125, output=-0.38071248114
			11'd1405: out = 32'b10000000000000000011000011011110; // input=-0.37255859375, output=-0.381764579591
			11'd1406: out = 32'b10000000000000000011000100000000; // input=-0.37353515625, output=-0.38281712261
			11'd1407: out = 32'b10000000000000000011000100100011; // input=-0.37451171875, output=-0.38387011193
			11'd1408: out = 32'b10000000000000000011000101000101; // input=-0.37548828125, output=-0.384923549288
			11'd1409: out = 32'b10000000000000000011000101101000; // input=-0.37646484375, output=-0.385977436426
			11'd1410: out = 32'b10000000000000000011000110001010; // input=-0.37744140625, output=-0.387031775094
			11'd1411: out = 32'b10000000000000000011000110101101; // input=-0.37841796875, output=-0.388086567045
			11'd1412: out = 32'b10000000000000000011000111001111; // input=-0.37939453125, output=-0.38914181404
			11'd1413: out = 32'b10000000000000000011000111110010; // input=-0.38037109375, output=-0.390197517845
			11'd1414: out = 32'b10000000000000000011001000010101; // input=-0.38134765625, output=-0.391253680232
			11'd1415: out = 32'b10000000000000000011001000110111; // input=-0.38232421875, output=-0.392310302978
			11'd1416: out = 32'b10000000000000000011001001011010; // input=-0.38330078125, output=-0.393367387867
			11'd1417: out = 32'b10000000000000000011001001111101; // input=-0.38427734375, output=-0.394424936689
			11'd1418: out = 32'b10000000000000000011001010011111; // input=-0.38525390625, output=-0.395482951241
			11'd1419: out = 32'b10000000000000000011001011000010; // input=-0.38623046875, output=-0.396541433322
			11'd1420: out = 32'b10000000000000000011001011100101; // input=-0.38720703125, output=-0.397600384742
			11'd1421: out = 32'b10000000000000000011001100000111; // input=-0.38818359375, output=-0.398659807314
			11'd1422: out = 32'b10000000000000000011001100101010; // input=-0.38916015625, output=-0.399719702858
			11'd1423: out = 32'b10000000000000000011001101001101; // input=-0.39013671875, output=-0.400780073201
			11'd1424: out = 32'b10000000000000000011001101110000; // input=-0.39111328125, output=-0.401840920174
			11'd1425: out = 32'b10000000000000000011001110010010; // input=-0.39208984375, output=-0.402902245618
			11'd1426: out = 32'b10000000000000000011001110110101; // input=-0.39306640625, output=-0.403964051377
			11'd1427: out = 32'b10000000000000000011001111011000; // input=-0.39404296875, output=-0.405026339302
			11'd1428: out = 32'b10000000000000000011001111111011; // input=-0.39501953125, output=-0.406089111252
			11'd1429: out = 32'b10000000000000000011010000011110; // input=-0.39599609375, output=-0.40715236909
			11'd1430: out = 32'b10000000000000000011010001000000; // input=-0.39697265625, output=-0.408216114687
			11'd1431: out = 32'b10000000000000000011010001100011; // input=-0.39794921875, output=-0.409280349921
			11'd1432: out = 32'b10000000000000000011010010000110; // input=-0.39892578125, output=-0.410345076676
			11'd1433: out = 32'b10000000000000000011010010101001; // input=-0.39990234375, output=-0.41141029684
			11'd1434: out = 32'b10000000000000000011010011001100; // input=-0.40087890625, output=-0.412476012313
			11'd1435: out = 32'b10000000000000000011010011101111; // input=-0.40185546875, output=-0.413542224997
			11'd1436: out = 32'b10000000000000000011010100010010; // input=-0.40283203125, output=-0.414608936802
			11'd1437: out = 32'b10000000000000000011010100110101; // input=-0.40380859375, output=-0.415676149646
			11'd1438: out = 32'b10000000000000000011010101011000; // input=-0.40478515625, output=-0.416743865453
			11'd1439: out = 32'b10000000000000000011010101111011; // input=-0.40576171875, output=-0.417812086153
			11'd1440: out = 32'b10000000000000000011010110011110; // input=-0.40673828125, output=-0.418880813684
			11'd1441: out = 32'b10000000000000000011010111000001; // input=-0.40771484375, output=-0.419950049991
			11'd1442: out = 32'b10000000000000000011010111100100; // input=-0.40869140625, output=-0.421019797024
			11'd1443: out = 32'b10000000000000000011011000000111; // input=-0.40966796875, output=-0.422090056743
			11'd1444: out = 32'b10000000000000000011011000101010; // input=-0.41064453125, output=-0.423160831114
			11'd1445: out = 32'b10000000000000000011011001001101; // input=-0.41162109375, output=-0.424232122107
			11'd1446: out = 32'b10000000000000000011011001110000; // input=-0.41259765625, output=-0.425303931704
			11'd1447: out = 32'b10000000000000000011011010010011; // input=-0.41357421875, output=-0.426376261892
			11'd1448: out = 32'b10000000000000000011011010110111; // input=-0.41455078125, output=-0.427449114664
			11'd1449: out = 32'b10000000000000000011011011011010; // input=-0.41552734375, output=-0.428522492022
			11'd1450: out = 32'b10000000000000000011011011111101; // input=-0.41650390625, output=-0.429596395974
			11'd1451: out = 32'b10000000000000000011011100100000; // input=-0.41748046875, output=-0.430670828538
			11'd1452: out = 32'b10000000000000000011011101000011; // input=-0.41845703125, output=-0.431745791736
			11'd1453: out = 32'b10000000000000000011011101100111; // input=-0.41943359375, output=-0.432821287599
			11'd1454: out = 32'b10000000000000000011011110001010; // input=-0.42041015625, output=-0.433897318166
			11'd1455: out = 32'b10000000000000000011011110101101; // input=-0.42138671875, output=-0.434973885483
			11'd1456: out = 32'b10000000000000000011011111010001; // input=-0.42236328125, output=-0.436050991604
			11'd1457: out = 32'b10000000000000000011011111110100; // input=-0.42333984375, output=-0.437128638589
			11'd1458: out = 32'b10000000000000000011100000010111; // input=-0.42431640625, output=-0.438206828509
			11'd1459: out = 32'b10000000000000000011100000111011; // input=-0.42529296875, output=-0.439285563439
			11'd1460: out = 32'b10000000000000000011100001011110; // input=-0.42626953125, output=-0.440364845464
			11'd1461: out = 32'b10000000000000000011100010000001; // input=-0.42724609375, output=-0.441444676676
			11'd1462: out = 32'b10000000000000000011100010100101; // input=-0.42822265625, output=-0.442525059177
			11'd1463: out = 32'b10000000000000000011100011001000; // input=-0.42919921875, output=-0.443605995073
			11'd1464: out = 32'b10000000000000000011100011101100; // input=-0.43017578125, output=-0.444687486481
			11'd1465: out = 32'b10000000000000000011100100001111; // input=-0.43115234375, output=-0.445769535526
			11'd1466: out = 32'b10000000000000000011100100110010; // input=-0.43212890625, output=-0.446852144339
			11'd1467: out = 32'b10000000000000000011100101010110; // input=-0.43310546875, output=-0.447935315062
			11'd1468: out = 32'b10000000000000000011100101111001; // input=-0.43408203125, output=-0.449019049842
			11'd1469: out = 32'b10000000000000000011100110011101; // input=-0.43505859375, output=-0.450103350837
			11'd1470: out = 32'b10000000000000000011100111000001; // input=-0.43603515625, output=-0.451188220212
			11'd1471: out = 32'b10000000000000000011100111100100; // input=-0.43701171875, output=-0.452273660141
			11'd1472: out = 32'b10000000000000000011101000001000; // input=-0.43798828125, output=-0.453359672806
			11'd1473: out = 32'b10000000000000000011101000101011; // input=-0.43896484375, output=-0.454446260396
			11'd1474: out = 32'b10000000000000000011101001001111; // input=-0.43994140625, output=-0.455533425112
			11'd1475: out = 32'b10000000000000000011101001110011; // input=-0.44091796875, output=-0.456621169161
			11'd1476: out = 32'b10000000000000000011101010010110; // input=-0.44189453125, output=-0.457709494758
			11'd1477: out = 32'b10000000000000000011101010111010; // input=-0.44287109375, output=-0.458798404129
			11'd1478: out = 32'b10000000000000000011101011011110; // input=-0.44384765625, output=-0.459887899507
			11'd1479: out = 32'b10000000000000000011101100000001; // input=-0.44482421875, output=-0.460977983136
			11'd1480: out = 32'b10000000000000000011101100100101; // input=-0.44580078125, output=-0.462068657266
			11'd1481: out = 32'b10000000000000000011101101001001; // input=-0.44677734375, output=-0.463159924156
			11'd1482: out = 32'b10000000000000000011101101101101; // input=-0.44775390625, output=-0.464251786078
			11'd1483: out = 32'b10000000000000000011101110010000; // input=-0.44873046875, output=-0.465344245308
			11'd1484: out = 32'b10000000000000000011101110110100; // input=-0.44970703125, output=-0.466437304135
			11'd1485: out = 32'b10000000000000000011101111011000; // input=-0.45068359375, output=-0.467530964854
			11'd1486: out = 32'b10000000000000000011101111111100; // input=-0.45166015625, output=-0.468625229772
			11'd1487: out = 32'b10000000000000000011110000100000; // input=-0.45263671875, output=-0.469720101202
			11'd1488: out = 32'b10000000000000000011110001000100; // input=-0.45361328125, output=-0.47081558147
			11'd1489: out = 32'b10000000000000000011110001101000; // input=-0.45458984375, output=-0.47191167291
			11'd1490: out = 32'b10000000000000000011110010001100; // input=-0.45556640625, output=-0.473008377863
			11'd1491: out = 32'b10000000000000000011110010101111; // input=-0.45654296875, output=-0.474105698684
			11'd1492: out = 32'b10000000000000000011110011010011; // input=-0.45751953125, output=-0.475203637734
			11'd1493: out = 32'b10000000000000000011110011110111; // input=-0.45849609375, output=-0.476302197385
			11'd1494: out = 32'b10000000000000000011110100011011; // input=-0.45947265625, output=-0.477401380019
			11'd1495: out = 32'b10000000000000000011110101000000; // input=-0.46044921875, output=-0.478501188027
			11'd1496: out = 32'b10000000000000000011110101100100; // input=-0.46142578125, output=-0.47960162381
			11'd1497: out = 32'b10000000000000000011110110001000; // input=-0.46240234375, output=-0.48070268978
			11'd1498: out = 32'b10000000000000000011110110101100; // input=-0.46337890625, output=-0.481804388357
			11'd1499: out = 32'b10000000000000000011110111010000; // input=-0.46435546875, output=-0.482906721972
			11'd1500: out = 32'b10000000000000000011110111110100; // input=-0.46533203125, output=-0.484009693068
			11'd1501: out = 32'b10000000000000000011111000011000; // input=-0.46630859375, output=-0.485113304095
			11'd1502: out = 32'b10000000000000000011111000111100; // input=-0.46728515625, output=-0.486217557514
			11'd1503: out = 32'b10000000000000000011111001100001; // input=-0.46826171875, output=-0.487322455798
			11'd1504: out = 32'b10000000000000000011111010000101; // input=-0.46923828125, output=-0.48842800143
			11'd1505: out = 32'b10000000000000000011111010101001; // input=-0.47021484375, output=-0.489534196901
			11'd1506: out = 32'b10000000000000000011111011001101; // input=-0.47119140625, output=-0.490641044716
			11'd1507: out = 32'b10000000000000000011111011110010; // input=-0.47216796875, output=-0.491748547388
			11'd1508: out = 32'b10000000000000000011111100010110; // input=-0.47314453125, output=-0.492856707441
			11'd1509: out = 32'b10000000000000000011111100111010; // input=-0.47412109375, output=-0.493965527411
			11'd1510: out = 32'b10000000000000000011111101011111; // input=-0.47509765625, output=-0.495075009844
			11'd1511: out = 32'b10000000000000000011111110000011; // input=-0.47607421875, output=-0.496185157297
			11'd1512: out = 32'b10000000000000000011111110100111; // input=-0.47705078125, output=-0.497295972337
			11'd1513: out = 32'b10000000000000000011111111001100; // input=-0.47802734375, output=-0.498407457545
			11'd1514: out = 32'b10000000000000000011111111110000; // input=-0.47900390625, output=-0.499519615509
			11'd1515: out = 32'b10000000000000000100000000010101; // input=-0.47998046875, output=-0.500632448832
			11'd1516: out = 32'b10000000000000000100000000111001; // input=-0.48095703125, output=-0.501745960124
			11'd1517: out = 32'b10000000000000000100000001011110; // input=-0.48193359375, output=-0.502860152012
			11'd1518: out = 32'b10000000000000000100000010000010; // input=-0.48291015625, output=-0.503975027128
			11'd1519: out = 32'b10000000000000000100000010100111; // input=-0.48388671875, output=-0.505090588121
			11'd1520: out = 32'b10000000000000000100000011001011; // input=-0.48486328125, output=-0.506206837649
			11'd1521: out = 32'b10000000000000000100000011110000; // input=-0.48583984375, output=-0.50732377838
			11'd1522: out = 32'b10000000000000000100000100010101; // input=-0.48681640625, output=-0.508441412998
			11'd1523: out = 32'b10000000000000000100000100111001; // input=-0.48779296875, output=-0.509559744196
			11'd1524: out = 32'b10000000000000000100000101011110; // input=-0.48876953125, output=-0.510678774679
			11'd1525: out = 32'b10000000000000000100000110000011; // input=-0.48974609375, output=-0.511798507164
			11'd1526: out = 32'b10000000000000000100000110100111; // input=-0.49072265625, output=-0.51291894438
			11'd1527: out = 32'b10000000000000000100000111001100; // input=-0.49169921875, output=-0.51404008907
			11'd1528: out = 32'b10000000000000000100000111110001; // input=-0.49267578125, output=-0.515161943987
			11'd1529: out = 32'b10000000000000000100001000010110; // input=-0.49365234375, output=-0.516284511897
			11'd1530: out = 32'b10000000000000000100001000111010; // input=-0.49462890625, output=-0.517407795578
			11'd1531: out = 32'b10000000000000000100001001011111; // input=-0.49560546875, output=-0.518531797822
			11'd1532: out = 32'b10000000000000000100001010000100; // input=-0.49658203125, output=-0.519656521432
			11'd1533: out = 32'b10000000000000000100001010101001; // input=-0.49755859375, output=-0.520781969224
			11'd1534: out = 32'b10000000000000000100001011001110; // input=-0.49853515625, output=-0.521908144027
			11'd1535: out = 32'b10000000000000000100001011110011; // input=-0.49951171875, output=-0.523035048684
			11'd1536: out = 32'b10000000000000000100001100011000; // input=-0.50048828125, output=-0.524162686048
			11'd1537: out = 32'b10000000000000000100001100111101; // input=-0.50146484375, output=-0.525291058987
			11'd1538: out = 32'b10000000000000000100001101100010; // input=-0.50244140625, output=-0.526420170383
			11'd1539: out = 32'b10000000000000000100001110000111; // input=-0.50341796875, output=-0.527550023129
			11'd1540: out = 32'b10000000000000000100001110101100; // input=-0.50439453125, output=-0.528680620133
			11'd1541: out = 32'b10000000000000000100001111010001; // input=-0.50537109375, output=-0.529811964315
			11'd1542: out = 32'b10000000000000000100001111110110; // input=-0.50634765625, output=-0.53094405861
			11'd1543: out = 32'b10000000000000000100010000011011; // input=-0.50732421875, output=-0.532076905965
			11'd1544: out = 32'b10000000000000000100010001000000; // input=-0.50830078125, output=-0.533210509343
			11'd1545: out = 32'b10000000000000000100010001100101; // input=-0.50927734375, output=-0.534344871718
			11'd1546: out = 32'b10000000000000000100010010001011; // input=-0.51025390625, output=-0.53547999608
			11'd1547: out = 32'b10000000000000000100010010110000; // input=-0.51123046875, output=-0.536615885432
			11'd1548: out = 32'b10000000000000000100010011010101; // input=-0.51220703125, output=-0.537752542791
			11'd1549: out = 32'b10000000000000000100010011111010; // input=-0.51318359375, output=-0.538889971188
			11'd1550: out = 32'b10000000000000000100010100100000; // input=-0.51416015625, output=-0.54002817367
			11'd1551: out = 32'b10000000000000000100010101000101; // input=-0.51513671875, output=-0.541167153296
			11'd1552: out = 32'b10000000000000000100010101101010; // input=-0.51611328125, output=-0.542306913141
			11'd1553: out = 32'b10000000000000000100010110010000; // input=-0.51708984375, output=-0.543447456295
			11'd1554: out = 32'b10000000000000000100010110110101; // input=-0.51806640625, output=-0.544588785861
			11'd1555: out = 32'b10000000000000000100010111011011; // input=-0.51904296875, output=-0.545730904958
			11'd1556: out = 32'b10000000000000000100011000000000; // input=-0.52001953125, output=-0.54687381672
			11'd1557: out = 32'b10000000000000000100011000100101; // input=-0.52099609375, output=-0.548017524295
			11'd1558: out = 32'b10000000000000000100011001001011; // input=-0.52197265625, output=-0.549162030848
			11'd1559: out = 32'b10000000000000000100011001110000; // input=-0.52294921875, output=-0.550307339557
			11'd1560: out = 32'b10000000000000000100011010010110; // input=-0.52392578125, output=-0.551453453618
			11'd1561: out = 32'b10000000000000000100011010111100; // input=-0.52490234375, output=-0.55260037624
			11'd1562: out = 32'b10000000000000000100011011100001; // input=-0.52587890625, output=-0.553748110648
			11'd1563: out = 32'b10000000000000000100011100000111; // input=-0.52685546875, output=-0.554896660084
			11'd1564: out = 32'b10000000000000000100011100101101; // input=-0.52783203125, output=-0.556046027806
			11'd1565: out = 32'b10000000000000000100011101010010; // input=-0.52880859375, output=-0.557196217085
			11'd1566: out = 32'b10000000000000000100011101111000; // input=-0.52978515625, output=-0.558347231212
			11'd1567: out = 32'b10000000000000000100011110011110; // input=-0.53076171875, output=-0.559499073492
			11'd1568: out = 32'b10000000000000000100011111000011; // input=-0.53173828125, output=-0.560651747246
			11'd1569: out = 32'b10000000000000000100011111101001; // input=-0.53271484375, output=-0.561805255813
			11'd1570: out = 32'b10000000000000000100100000001111; // input=-0.53369140625, output=-0.562959602546
			11'd1571: out = 32'b10000000000000000100100000110101; // input=-0.53466796875, output=-0.564114790818
			11'd1572: out = 32'b10000000000000000100100001011011; // input=-0.53564453125, output=-0.565270824016
			11'd1573: out = 32'b10000000000000000100100010000001; // input=-0.53662109375, output=-0.566427705546
			11'd1574: out = 32'b10000000000000000100100010100111; // input=-0.53759765625, output=-0.567585438829
			11'd1575: out = 32'b10000000000000000100100011001101; // input=-0.53857421875, output=-0.568744027306
			11'd1576: out = 32'b10000000000000000100100011110011; // input=-0.53955078125, output=-0.569903474432
			11'd1577: out = 32'b10000000000000000100100100011001; // input=-0.54052734375, output=-0.571063783681
			11'd1578: out = 32'b10000000000000000100100100111111; // input=-0.54150390625, output=-0.572224958546
			11'd1579: out = 32'b10000000000000000100100101100101; // input=-0.54248046875, output=-0.573387002535
			11'd1580: out = 32'b10000000000000000100100110001011; // input=-0.54345703125, output=-0.574549919176
			11'd1581: out = 32'b10000000000000000100100110110001; // input=-0.54443359375, output=-0.575713712013
			11'd1582: out = 32'b10000000000000000100100111010111; // input=-0.54541015625, output=-0.576878384612
			11'd1583: out = 32'b10000000000000000100100111111101; // input=-0.54638671875, output=-0.578043940552
			11'd1584: out = 32'b10000000000000000100101000100100; // input=-0.54736328125, output=-0.579210383434
			11'd1585: out = 32'b10000000000000000100101001001010; // input=-0.54833984375, output=-0.580377716876
			11'd1586: out = 32'b10000000000000000100101001110000; // input=-0.54931640625, output=-0.581545944516
			11'd1587: out = 32'b10000000000000000100101010010110; // input=-0.55029296875, output=-0.58271507001
			11'd1588: out = 32'b10000000000000000100101010111101; // input=-0.55126953125, output=-0.583885097033
			11'd1589: out = 32'b10000000000000000100101011100011; // input=-0.55224609375, output=-0.585056029278
			11'd1590: out = 32'b10000000000000000100101100001010; // input=-0.55322265625, output=-0.586227870461
			11'd1591: out = 32'b10000000000000000100101100110000; // input=-0.55419921875, output=-0.587400624313
			11'd1592: out = 32'b10000000000000000100101101010110; // input=-0.55517578125, output=-0.588574294586
			11'd1593: out = 32'b10000000000000000100101101111101; // input=-0.55615234375, output=-0.589748885055
			11'd1594: out = 32'b10000000000000000100101110100011; // input=-0.55712890625, output=-0.590924399509
			11'd1595: out = 32'b10000000000000000100101111001010; // input=-0.55810546875, output=-0.592100841762
			11'd1596: out = 32'b10000000000000000100101111110001; // input=-0.55908203125, output=-0.593278215646
			11'd1597: out = 32'b10000000000000000100110000010111; // input=-0.56005859375, output=-0.594456525014
			11'd1598: out = 32'b10000000000000000100110000111110; // input=-0.56103515625, output=-0.595635773739
			11'd1599: out = 32'b10000000000000000100110001100100; // input=-0.56201171875, output=-0.596815965716
			11'd1600: out = 32'b10000000000000000100110010001011; // input=-0.56298828125, output=-0.597997104858
			11'd1601: out = 32'b10000000000000000100110010110010; // input=-0.56396484375, output=-0.599179195102
			11'd1602: out = 32'b10000000000000000100110011011001; // input=-0.56494140625, output=-0.600362240405
			11'd1603: out = 32'b10000000000000000100110011111111; // input=-0.56591796875, output=-0.601546244745
			11'd1604: out = 32'b10000000000000000100110100100110; // input=-0.56689453125, output=-0.602731212123
			11'd1605: out = 32'b10000000000000000100110101001101; // input=-0.56787109375, output=-0.60391714656
			11'd1606: out = 32'b10000000000000000100110101110100; // input=-0.56884765625, output=-0.6051040521
			11'd1607: out = 32'b10000000000000000100110110011011; // input=-0.56982421875, output=-0.606291932808
			11'd1608: out = 32'b10000000000000000100110111000010; // input=-0.57080078125, output=-0.607480792772
			11'd1609: out = 32'b10000000000000000100110111101001; // input=-0.57177734375, output=-0.608670636103
			11'd1610: out = 32'b10000000000000000100111000010000; // input=-0.57275390625, output=-0.609861466933
			11'd1611: out = 32'b10000000000000000100111000110111; // input=-0.57373046875, output=-0.611053289418
			11'd1612: out = 32'b10000000000000000100111001011110; // input=-0.57470703125, output=-0.612246107738
			11'd1613: out = 32'b10000000000000000100111010000101; // input=-0.57568359375, output=-0.613439926093
			11'd1614: out = 32'b10000000000000000100111010101100; // input=-0.57666015625, output=-0.614634748708
			11'd1615: out = 32'b10000000000000000100111011010100; // input=-0.57763671875, output=-0.615830579834
			11'd1616: out = 32'b10000000000000000100111011111011; // input=-0.57861328125, output=-0.617027423741
			11'd1617: out = 32'b10000000000000000100111100100010; // input=-0.57958984375, output=-0.618225284727
			11'd1618: out = 32'b10000000000000000100111101001001; // input=-0.58056640625, output=-0.619424167112
			11'd1619: out = 32'b10000000000000000100111101110001; // input=-0.58154296875, output=-0.62062407524
			11'd1620: out = 32'b10000000000000000100111110011000; // input=-0.58251953125, output=-0.621825013482
			11'd1621: out = 32'b10000000000000000100111110111111; // input=-0.58349609375, output=-0.623026986232
			11'd1622: out = 32'b10000000000000000100111111100111; // input=-0.58447265625, output=-0.624229997907
			11'd1623: out = 32'b10000000000000000101000000001110; // input=-0.58544921875, output=-0.625434052954
			11'd1624: out = 32'b10000000000000000101000000110110; // input=-0.58642578125, output=-0.62663915584
			11'd1625: out = 32'b10000000000000000101000001011101; // input=-0.58740234375, output=-0.627845311062
			11'd1626: out = 32'b10000000000000000101000010000101; // input=-0.58837890625, output=-0.629052523141
			11'd1627: out = 32'b10000000000000000101000010101100; // input=-0.58935546875, output=-0.630260796623
			11'd1628: out = 32'b10000000000000000101000011010100; // input=-0.59033203125, output=-0.631470136082
			11'd1629: out = 32'b10000000000000000101000011111100; // input=-0.59130859375, output=-0.632680546116
			11'd1630: out = 32'b10000000000000000101000100100011; // input=-0.59228515625, output=-0.633892031354
			11'd1631: out = 32'b10000000000000000101000101001011; // input=-0.59326171875, output=-0.635104596447
			11'd1632: out = 32'b10000000000000000101000101110011; // input=-0.59423828125, output=-0.636318246077
			11'd1633: out = 32'b10000000000000000101000110011011; // input=-0.59521484375, output=-0.63753298495
			11'd1634: out = 32'b10000000000000000101000111000011; // input=-0.59619140625, output=-0.638748817803
			11'd1635: out = 32'b10000000000000000101000111101010; // input=-0.59716796875, output=-0.639965749399
			11'd1636: out = 32'b10000000000000000101001000010010; // input=-0.59814453125, output=-0.641183784528
			11'd1637: out = 32'b10000000000000000101001000111010; // input=-0.59912109375, output=-0.64240292801
			11'd1638: out = 32'b10000000000000000101001001100010; // input=-0.60009765625, output=-0.643623184695
			11'd1639: out = 32'b10000000000000000101001010001010; // input=-0.60107421875, output=-0.644844559457
			11'd1640: out = 32'b10000000000000000101001010110010; // input=-0.60205078125, output=-0.646067057204
			11'd1641: out = 32'b10000000000000000101001011011010; // input=-0.60302734375, output=-0.647290682871
			11'd1642: out = 32'b10000000000000000101001100000011; // input=-0.60400390625, output=-0.648515441423
			11'd1643: out = 32'b10000000000000000101001100101011; // input=-0.60498046875, output=-0.649741337855
			11'd1644: out = 32'b10000000000000000101001101010011; // input=-0.60595703125, output=-0.650968377191
			11'd1645: out = 32'b10000000000000000101001101111011; // input=-0.60693359375, output=-0.652196564486
			11'd1646: out = 32'b10000000000000000101001110100011; // input=-0.60791015625, output=-0.653425904828
			11'd1647: out = 32'b10000000000000000101001111001100; // input=-0.60888671875, output=-0.654656403331
			11'd1648: out = 32'b10000000000000000101001111110100; // input=-0.60986328125, output=-0.655888065144
			11'd1649: out = 32'b10000000000000000101010000011101; // input=-0.61083984375, output=-0.657120895447
			11'd1650: out = 32'b10000000000000000101010001000101; // input=-0.61181640625, output=-0.658354899451
			11'd1651: out = 32'b10000000000000000101010001101101; // input=-0.61279296875, output=-0.659590082398
			11'd1652: out = 32'b10000000000000000101010010010110; // input=-0.61376953125, output=-0.660826449565
			11'd1653: out = 32'b10000000000000000101010010111111; // input=-0.61474609375, output=-0.662064006259
			11'd1654: out = 32'b10000000000000000101010011100111; // input=-0.61572265625, output=-0.66330275782
			11'd1655: out = 32'b10000000000000000101010100010000; // input=-0.61669921875, output=-0.664542709624
			11'd1656: out = 32'b10000000000000000101010100111000; // input=-0.61767578125, output=-0.665783867077
			11'd1657: out = 32'b10000000000000000101010101100001; // input=-0.61865234375, output=-0.667026235621
			11'd1658: out = 32'b10000000000000000101010110001010; // input=-0.61962890625, output=-0.668269820732
			11'd1659: out = 32'b10000000000000000101010110110011; // input=-0.62060546875, output=-0.669514627918
			11'd1660: out = 32'b10000000000000000101010111011011; // input=-0.62158203125, output=-0.670760662725
			11'd1661: out = 32'b10000000000000000101011000000100; // input=-0.62255859375, output=-0.672007930733
			11'd1662: out = 32'b10000000000000000101011000101101; // input=-0.62353515625, output=-0.673256437555
			11'd1663: out = 32'b10000000000000000101011001010110; // input=-0.62451171875, output=-0.674506188843
			11'd1664: out = 32'b10000000000000000101011001111111; // input=-0.62548828125, output=-0.675757190283
			11'd1665: out = 32'b10000000000000000101011010101000; // input=-0.62646484375, output=-0.677009447598
			11'd1666: out = 32'b10000000000000000101011011010001; // input=-0.62744140625, output=-0.678262966548
			11'd1667: out = 32'b10000000000000000101011011111010; // input=-0.62841796875, output=-0.679517752929
			11'd1668: out = 32'b10000000000000000101011100100100; // input=-0.62939453125, output=-0.680773812575
			11'd1669: out = 32'b10000000000000000101011101001101; // input=-0.63037109375, output=-0.682031151358
			11'd1670: out = 32'b10000000000000000101011101110110; // input=-0.63134765625, output=-0.683289775188
			11'd1671: out = 32'b10000000000000000101011110011111; // input=-0.63232421875, output=-0.684549690012
			11'd1672: out = 32'b10000000000000000101011111001001; // input=-0.63330078125, output=-0.685810901818
			11'd1673: out = 32'b10000000000000000101011111110010; // input=-0.63427734375, output=-0.687073416632
			11'd1674: out = 32'b10000000000000000101100000011011; // input=-0.63525390625, output=-0.688337240519
			11'd1675: out = 32'b10000000000000000101100001000101; // input=-0.63623046875, output=-0.689602379584
			11'd1676: out = 32'b10000000000000000101100001101110; // input=-0.63720703125, output=-0.690868839974
			11'd1677: out = 32'b10000000000000000101100010011000; // input=-0.63818359375, output=-0.692136627875
			11'd1678: out = 32'b10000000000000000101100011000010; // input=-0.63916015625, output=-0.693405749514
			11'd1679: out = 32'b10000000000000000101100011101011; // input=-0.64013671875, output=-0.694676211161
			11'd1680: out = 32'b10000000000000000101100100010101; // input=-0.64111328125, output=-0.695948019125
			11'd1681: out = 32'b10000000000000000101100100111111; // input=-0.64208984375, output=-0.697221179759
			11'd1682: out = 32'b10000000000000000101100101101000; // input=-0.64306640625, output=-0.69849569946
			11'd1683: out = 32'b10000000000000000101100110010010; // input=-0.64404296875, output=-0.699771584666
			11'd1684: out = 32'b10000000000000000101100110111100; // input=-0.64501953125, output=-0.701048841859
			11'd1685: out = 32'b10000000000000000101100111100110; // input=-0.64599609375, output=-0.702327477564
			11'd1686: out = 32'b10000000000000000101101000010000; // input=-0.64697265625, output=-0.703607498353
			11'd1687: out = 32'b10000000000000000101101000111010; // input=-0.64794921875, output=-0.70488891084
			11'd1688: out = 32'b10000000000000000101101001100100; // input=-0.64892578125, output=-0.706171721686
			11'd1689: out = 32'b10000000000000000101101010001110; // input=-0.64990234375, output=-0.707455937596
			11'd1690: out = 32'b10000000000000000101101010111000; // input=-0.65087890625, output=-0.708741565323
			11'd1691: out = 32'b10000000000000000101101011100010; // input=-0.65185546875, output=-0.710028611664
			11'd1692: out = 32'b10000000000000000101101100001100; // input=-0.65283203125, output=-0.711317083466
			11'd1693: out = 32'b10000000000000000101101100110111; // input=-0.65380859375, output=-0.712606987621
			11'd1694: out = 32'b10000000000000000101101101100001; // input=-0.65478515625, output=-0.713898331071
			11'd1695: out = 32'b10000000000000000101101110001011; // input=-0.65576171875, output=-0.715191120804
			11'd1696: out = 32'b10000000000000000101101110110110; // input=-0.65673828125, output=-0.71648536386
			11'd1697: out = 32'b10000000000000000101101111100000; // input=-0.65771484375, output=-0.717781067325
			11'd1698: out = 32'b10000000000000000101110000001011; // input=-0.65869140625, output=-0.719078238338
			11'd1699: out = 32'b10000000000000000101110000110101; // input=-0.65966796875, output=-0.720376884086
			11'd1700: out = 32'b10000000000000000101110001100000; // input=-0.66064453125, output=-0.721677011809
			11'd1701: out = 32'b10000000000000000101110010001011; // input=-0.66162109375, output=-0.722978628796
			11'd1702: out = 32'b10000000000000000101110010110101; // input=-0.66259765625, output=-0.72428174239
			11'd1703: out = 32'b10000000000000000101110011100000; // input=-0.66357421875, output=-0.725586359986
			11'd1704: out = 32'b10000000000000000101110100001011; // input=-0.66455078125, output=-0.726892489032
			11'd1705: out = 32'b10000000000000000101110100110110; // input=-0.66552734375, output=-0.728200137029
			11'd1706: out = 32'b10000000000000000101110101100001; // input=-0.66650390625, output=-0.729509311532
			11'd1707: out = 32'b10000000000000000101110110001100; // input=-0.66748046875, output=-0.730820020153
			11'd1708: out = 32'b10000000000000000101110110110111; // input=-0.66845703125, output=-0.732132270556
			11'd1709: out = 32'b10000000000000000101110111100010; // input=-0.66943359375, output=-0.733446070462
			11'd1710: out = 32'b10000000000000000101111000001101; // input=-0.67041015625, output=-0.734761427651
			11'd1711: out = 32'b10000000000000000101111000111000; // input=-0.67138671875, output=-0.736078349955
			11'd1712: out = 32'b10000000000000000101111001100011; // input=-0.67236328125, output=-0.737396845268
			11'd1713: out = 32'b10000000000000000101111010001110; // input=-0.67333984375, output=-0.73871692154
			11'd1714: out = 32'b10000000000000000101111010111010; // input=-0.67431640625, output=-0.74003858678
			11'd1715: out = 32'b10000000000000000101111011100101; // input=-0.67529296875, output=-0.741361849058
			11'd1716: out = 32'b10000000000000000101111100010000; // input=-0.67626953125, output=-0.742686716502
			11'd1717: out = 32'b10000000000000000101111100111100; // input=-0.67724609375, output=-0.744013197301
			11'd1718: out = 32'b10000000000000000101111101100111; // input=-0.67822265625, output=-0.745341299708
			11'd1719: out = 32'b10000000000000000101111110010011; // input=-0.67919921875, output=-0.746671032034
			11'd1720: out = 32'b10000000000000000101111110111111; // input=-0.68017578125, output=-0.748002402655
			11'd1721: out = 32'b10000000000000000101111111101010; // input=-0.68115234375, output=-0.749335420011
			11'd1722: out = 32'b10000000000000000110000000010110; // input=-0.68212890625, output=-0.750670092604
			11'd1723: out = 32'b10000000000000000110000001000010; // input=-0.68310546875, output=-0.752006429003
			11'd1724: out = 32'b10000000000000000110000001101110; // input=-0.68408203125, output=-0.75334443784
			11'd1725: out = 32'b10000000000000000110000010011001; // input=-0.68505859375, output=-0.754684127815
			11'd1726: out = 32'b10000000000000000110000011000101; // input=-0.68603515625, output=-0.756025507694
			11'd1727: out = 32'b10000000000000000110000011110001; // input=-0.68701171875, output=-0.757368586311
			11'd1728: out = 32'b10000000000000000110000100011110; // input=-0.68798828125, output=-0.758713372569
			11'd1729: out = 32'b10000000000000000110000101001010; // input=-0.68896484375, output=-0.760059875439
			11'd1730: out = 32'b10000000000000000110000101110110; // input=-0.68994140625, output=-0.761408103962
			11'd1731: out = 32'b10000000000000000110000110100010; // input=-0.69091796875, output=-0.76275806725
			11'd1732: out = 32'b10000000000000000110000111001110; // input=-0.69189453125, output=-0.764109774486
			11'd1733: out = 32'b10000000000000000110000111111011; // input=-0.69287109375, output=-0.765463234926
			11'd1734: out = 32'b10000000000000000110001000100111; // input=-0.69384765625, output=-0.766818457899
			11'd1735: out = 32'b10000000000000000110001001010100; // input=-0.69482421875, output=-0.768175452807
			11'd1736: out = 32'b10000000000000000110001010000000; // input=-0.69580078125, output=-0.769534229128
			11'd1737: out = 32'b10000000000000000110001010101101; // input=-0.69677734375, output=-0.770894796414
			11'd1738: out = 32'b10000000000000000110001011011001; // input=-0.69775390625, output=-0.772257164294
			11'd1739: out = 32'b10000000000000000110001100000110; // input=-0.69873046875, output=-0.773621342475
			11'd1740: out = 32'b10000000000000000110001100110011; // input=-0.69970703125, output=-0.774987340742
			11'd1741: out = 32'b10000000000000000110001101100000; // input=-0.70068359375, output=-0.776355168958
			11'd1742: out = 32'b10000000000000000110001110001100; // input=-0.70166015625, output=-0.777724837066
			11'd1743: out = 32'b10000000000000000110001110111001; // input=-0.70263671875, output=-0.779096355093
			11'd1744: out = 32'b10000000000000000110001111100110; // input=-0.70361328125, output=-0.780469733143
			11'd1745: out = 32'b10000000000000000110010000010011; // input=-0.70458984375, output=-0.781844981407
			11'd1746: out = 32'b10000000000000000110010001000001; // input=-0.70556640625, output=-0.783222110157
			11'd1747: out = 32'b10000000000000000110010001101110; // input=-0.70654296875, output=-0.78460112975
			11'd1748: out = 32'b10000000000000000110010010011011; // input=-0.70751953125, output=-0.78598205063
			11'd1749: out = 32'b10000000000000000110010011001000; // input=-0.70849609375, output=-0.787364883328
			11'd1750: out = 32'b10000000000000000110010011110110; // input=-0.70947265625, output=-0.788749638461
			11'd1751: out = 32'b10000000000000000110010100100011; // input=-0.71044921875, output=-0.790136326735
			11'd1752: out = 32'b10000000000000000110010101010001; // input=-0.71142578125, output=-0.791524958947
			11'd1753: out = 32'b10000000000000000110010101111110; // input=-0.71240234375, output=-0.792915545985
			11'd1754: out = 32'b10000000000000000110010110101100; // input=-0.71337890625, output=-0.794308098827
			11'd1755: out = 32'b10000000000000000110010111011010; // input=-0.71435546875, output=-0.795702628547
			11'd1756: out = 32'b10000000000000000110011000000111; // input=-0.71533203125, output=-0.797099146312
			11'd1757: out = 32'b10000000000000000110011000110101; // input=-0.71630859375, output=-0.798497663382
			11'd1758: out = 32'b10000000000000000110011001100011; // input=-0.71728515625, output=-0.799898191117
			11'd1759: out = 32'b10000000000000000110011010010001; // input=-0.71826171875, output=-0.801300740973
			11'd1760: out = 32'b10000000000000000110011010111111; // input=-0.71923828125, output=-0.802705324505
			11'd1761: out = 32'b10000000000000000110011011101101; // input=-0.72021484375, output=-0.804111953369
			11'd1762: out = 32'b10000000000000000110011100011011; // input=-0.72119140625, output=-0.805520639322
			11'd1763: out = 32'b10000000000000000110011101001010; // input=-0.72216796875, output=-0.806931394221
			11'd1764: out = 32'b10000000000000000110011101111000; // input=-0.72314453125, output=-0.808344230032
			11'd1765: out = 32'b10000000000000000110011110100110; // input=-0.72412109375, output=-0.809759158821
			11'd1766: out = 32'b10000000000000000110011111010101; // input=-0.72509765625, output=-0.811176192763
			11'd1767: out = 32'b10000000000000000110100000000011; // input=-0.72607421875, output=-0.812595344141
			11'd1768: out = 32'b10000000000000000110100000110010; // input=-0.72705078125, output=-0.814016625347
			11'd1769: out = 32'b10000000000000000110100001100000; // input=-0.72802734375, output=-0.815440048882
			11'd1770: out = 32'b10000000000000000110100010001111; // input=-0.72900390625, output=-0.816865627361
			11'd1771: out = 32'b10000000000000000110100010111110; // input=-0.72998046875, output=-0.81829337351
			11'd1772: out = 32'b10000000000000000110100011101101; // input=-0.73095703125, output=-0.819723300173
			11'd1773: out = 32'b10000000000000000110100100011100; // input=-0.73193359375, output=-0.821155420307
			11'd1774: out = 32'b10000000000000000110100101001011; // input=-0.73291015625, output=-0.822589746989
			11'd1775: out = 32'b10000000000000000110100101111010; // input=-0.73388671875, output=-0.824026293413
			11'd1776: out = 32'b10000000000000000110100110101001; // input=-0.73486328125, output=-0.825465072897
			11'd1777: out = 32'b10000000000000000110100111011000; // input=-0.73583984375, output=-0.826906098877
			11'd1778: out = 32'b10000000000000000110101000000111; // input=-0.73681640625, output=-0.828349384918
			11'd1779: out = 32'b10000000000000000110101000110111; // input=-0.73779296875, output=-0.829794944707
			11'd1780: out = 32'b10000000000000000110101001100110; // input=-0.73876953125, output=-0.831242792059
			11'd1781: out = 32'b10000000000000000110101010010110; // input=-0.73974609375, output=-0.832692940918
			11'd1782: out = 32'b10000000000000000110101011000101; // input=-0.74072265625, output=-0.834145405359
			11'd1783: out = 32'b10000000000000000110101011110101; // input=-0.74169921875, output=-0.835600199588
			11'd1784: out = 32'b10000000000000000110101100100101; // input=-0.74267578125, output=-0.837057337948
			11'd1785: out = 32'b10000000000000000110101101010101; // input=-0.74365234375, output=-0.838516834915
			11'd1786: out = 32'b10000000000000000110101110000100; // input=-0.74462890625, output=-0.839978705103
			11'd1787: out = 32'b10000000000000000110101110110100; // input=-0.74560546875, output=-0.841442963267
			11'd1788: out = 32'b10000000000000000110101111100100; // input=-0.74658203125, output=-0.842909624303
			11'd1789: out = 32'b10000000000000000110110000010101; // input=-0.74755859375, output=-0.844378703249
			11'd1790: out = 32'b10000000000000000110110001000101; // input=-0.74853515625, output=-0.845850215289
			11'd1791: out = 32'b10000000000000000110110001110101; // input=-0.74951171875, output=-0.847324175756
			11'd1792: out = 32'b10000000000000000110110010100101; // input=-0.75048828125, output=-0.84880060013
			11'd1793: out = 32'b10000000000000000110110011010110; // input=-0.75146484375, output=-0.850279504044
			11'd1794: out = 32'b10000000000000000110110100000111; // input=-0.75244140625, output=-0.851760903282
			11'd1795: out = 32'b10000000000000000110110100110111; // input=-0.75341796875, output=-0.853244813787
			11'd1796: out = 32'b10000000000000000110110101101000; // input=-0.75439453125, output=-0.854731251657
			11'd1797: out = 32'b10000000000000000110110110011001; // input=-0.75537109375, output=-0.856220233152
			11'd1798: out = 32'b10000000000000000110110111001001; // input=-0.75634765625, output=-0.857711774692
			11'd1799: out = 32'b10000000000000000110110111111010; // input=-0.75732421875, output=-0.859205892863
			11'd1800: out = 32'b10000000000000000110111000101100; // input=-0.75830078125, output=-0.860702604419
			11'd1801: out = 32'b10000000000000000110111001011101; // input=-0.75927734375, output=-0.86220192628
			11'd1802: out = 32'b10000000000000000110111010001110; // input=-0.76025390625, output=-0.863703875539
			11'd1803: out = 32'b10000000000000000110111010111111; // input=-0.76123046875, output=-0.865208469465
			11'd1804: out = 32'b10000000000000000110111011110001; // input=-0.76220703125, output=-0.866715725501
			11'd1805: out = 32'b10000000000000000110111100100010; // input=-0.76318359375, output=-0.868225661271
			11'd1806: out = 32'b10000000000000000110111101010100; // input=-0.76416015625, output=-0.869738294579
			11'd1807: out = 32'b10000000000000000110111110000101; // input=-0.76513671875, output=-0.871253643414
			11'd1808: out = 32'b10000000000000000110111110110111; // input=-0.76611328125, output=-0.872771725953
			11'd1809: out = 32'b10000000000000000110111111101001; // input=-0.76708984375, output=-0.874292560562
			11'd1810: out = 32'b10000000000000000111000000011011; // input=-0.76806640625, output=-0.875816165799
			11'd1811: out = 32'b10000000000000000111000001001101; // input=-0.76904296875, output=-0.877342560418
			11'd1812: out = 32'b10000000000000000111000001111111; // input=-0.77001953125, output=-0.878871763373
			11'd1813: out = 32'b10000000000000000111000010110001; // input=-0.77099609375, output=-0.880403793817
			11'd1814: out = 32'b10000000000000000111000011100011; // input=-0.77197265625, output=-0.881938671108
			11'd1815: out = 32'b10000000000000000111000100010110; // input=-0.77294921875, output=-0.883476414811
			11'd1816: out = 32'b10000000000000000111000101001000; // input=-0.77392578125, output=-0.885017044704
			11'd1817: out = 32'b10000000000000000111000101111011; // input=-0.77490234375, output=-0.886560580776
			11'd1818: out = 32'b10000000000000000111000110101101; // input=-0.77587890625, output=-0.888107043235
			11'd1819: out = 32'b10000000000000000111000111100000; // input=-0.77685546875, output=-0.889656452506
			11'd1820: out = 32'b10000000000000000111001000010011; // input=-0.77783203125, output=-0.891208829243
			11'd1821: out = 32'b10000000000000000111001001000110; // input=-0.77880859375, output=-0.892764194322
			11'd1822: out = 32'b10000000000000000111001001111001; // input=-0.77978515625, output=-0.894322568854
			11'd1823: out = 32'b10000000000000000111001010101100; // input=-0.78076171875, output=-0.895883974181
			11'd1824: out = 32'b10000000000000000111001011100000; // input=-0.78173828125, output=-0.897448431885
			11'd1825: out = 32'b10000000000000000111001100010011; // input=-0.78271484375, output=-0.899015963789
			11'd1826: out = 32'b10000000000000000111001101000110; // input=-0.78369140625, output=-0.900586591962
			11'd1827: out = 32'b10000000000000000111001101111010; // input=-0.78466796875, output=-0.902160338722
			11'd1828: out = 32'b10000000000000000111001110101110; // input=-0.78564453125, output=-0.903737226641
			11'd1829: out = 32'b10000000000000000111001111100001; // input=-0.78662109375, output=-0.905317278548
			11'd1830: out = 32'b10000000000000000111010000010101; // input=-0.78759765625, output=-0.906900517533
			11'd1831: out = 32'b10000000000000000111010001001001; // input=-0.78857421875, output=-0.908486966953
			11'd1832: out = 32'b10000000000000000111010001111101; // input=-0.78955078125, output=-0.910076650436
			11'd1833: out = 32'b10000000000000000111010010110010; // input=-0.79052734375, output=-0.911669591883
			11'd1834: out = 32'b10000000000000000111010011100110; // input=-0.79150390625, output=-0.913265815473
			11'd1835: out = 32'b10000000000000000111010100011010; // input=-0.79248046875, output=-0.914865345673
			11'd1836: out = 32'b10000000000000000111010101001111; // input=-0.79345703125, output=-0.916468207233
			11'd1837: out = 32'b10000000000000000111010110000011; // input=-0.79443359375, output=-0.918074425201
			11'd1838: out = 32'b10000000000000000111010110111000; // input=-0.79541015625, output=-0.919684024919
			11'd1839: out = 32'b10000000000000000111010111101101; // input=-0.79638671875, output=-0.921297032036
			11'd1840: out = 32'b10000000000000000111011000100010; // input=-0.79736328125, output=-0.922913472506
			11'd1841: out = 32'b10000000000000000111011001010111; // input=-0.79833984375, output=-0.924533372597
			11'd1842: out = 32'b10000000000000000111011010001100; // input=-0.79931640625, output=-0.926156758898
			11'd1843: out = 32'b10000000000000000111011011000010; // input=-0.80029296875, output=-0.92778365832
			11'd1844: out = 32'b10000000000000000111011011110111; // input=-0.80126953125, output=-0.929414098105
			11'd1845: out = 32'b10000000000000000111011100101101; // input=-0.80224609375, output=-0.931048105828
			11'd1846: out = 32'b10000000000000000111011101100010; // input=-0.80322265625, output=-0.932685709409
			11'd1847: out = 32'b10000000000000000111011110011000; // input=-0.80419921875, output=-0.934326937112
			11'd1848: out = 32'b10000000000000000111011111001110; // input=-0.80517578125, output=-0.935971817557
			11'd1849: out = 32'b10000000000000000111100000000100; // input=-0.80615234375, output=-0.937620379721
			11'd1850: out = 32'b10000000000000000111100000111010; // input=-0.80712890625, output=-0.93927265295
			11'd1851: out = 32'b10000000000000000111100001110000; // input=-0.80810546875, output=-0.940928666959
			11'd1852: out = 32'b10000000000000000111100010100111; // input=-0.80908203125, output=-0.942588451845
			11'd1853: out = 32'b10000000000000000111100011011101; // input=-0.81005859375, output=-0.944252038088
			11'd1854: out = 32'b10000000000000000111100100010100; // input=-0.81103515625, output=-0.945919456565
			11'd1855: out = 32'b10000000000000000111100101001011; // input=-0.81201171875, output=-0.947590738548
			11'd1856: out = 32'b10000000000000000111100110000010; // input=-0.81298828125, output=-0.949265915721
			11'd1857: out = 32'b10000000000000000111100110111001; // input=-0.81396484375, output=-0.95094502018
			11'd1858: out = 32'b10000000000000000111100111110000; // input=-0.81494140625, output=-0.952628084445
			11'd1859: out = 32'b10000000000000000111101000100111; // input=-0.81591796875, output=-0.954315141464
			11'd1860: out = 32'b10000000000000000111101001011110; // input=-0.81689453125, output=-0.956006224626
			11'd1861: out = 32'b10000000000000000111101010010110; // input=-0.81787109375, output=-0.957701367765
			11'd1862: out = 32'b10000000000000000111101011001110; // input=-0.81884765625, output=-0.95940060517
			11'd1863: out = 32'b10000000000000000111101100000101; // input=-0.81982421875, output=-0.961103971595
			11'd1864: out = 32'b10000000000000000111101100111101; // input=-0.82080078125, output=-0.962811502264
			11'd1865: out = 32'b10000000000000000111101101110101; // input=-0.82177734375, output=-0.964523232885
			11'd1866: out = 32'b10000000000000000111101110101110; // input=-0.82275390625, output=-0.966239199654
			11'd1867: out = 32'b10000000000000000111101111100110; // input=-0.82373046875, output=-0.967959439271
			11'd1868: out = 32'b10000000000000000111110000011111; // input=-0.82470703125, output=-0.969683988941
			11'd1869: out = 32'b10000000000000000111110001010111; // input=-0.82568359375, output=-0.971412886393
			11'd1870: out = 32'b10000000000000000111110010010000; // input=-0.82666015625, output=-0.973146169884
			11'd1871: out = 32'b10000000000000000111110011001001; // input=-0.82763671875, output=-0.974883878213
			11'd1872: out = 32'b10000000000000000111110100000010; // input=-0.82861328125, output=-0.976626050731
			11'd1873: out = 32'b10000000000000000111110100111011; // input=-0.82958984375, output=-0.978372727348
			11'd1874: out = 32'b10000000000000000111110101110101; // input=-0.83056640625, output=-0.980123948551
			11'd1875: out = 32'b10000000000000000111110110101110; // input=-0.83154296875, output=-0.981879755413
			11'd1876: out = 32'b10000000000000000111110111101000; // input=-0.83251953125, output=-0.983640189601
			11'd1877: out = 32'b10000000000000000111111000100010; // input=-0.83349609375, output=-0.985405293394
			11'd1878: out = 32'b10000000000000000111111001011100; // input=-0.83447265625, output=-0.987175109694
			11'd1879: out = 32'b10000000000000000111111010010110; // input=-0.83544921875, output=-0.988949682035
			11'd1880: out = 32'b10000000000000000111111011010000; // input=-0.83642578125, output=-0.990729054601
			11'd1881: out = 32'b10000000000000000111111100001011; // input=-0.83740234375, output=-0.992513272239
			11'd1882: out = 32'b10000000000000000111111101000101; // input=-0.83837890625, output=-0.99430238047
			11'd1883: out = 32'b10000000000000000111111110000000; // input=-0.83935546875, output=-0.996096425507
			11'd1884: out = 32'b10000000000000000111111110111011; // input=-0.84033203125, output=-0.997895454266
			11'd1885: out = 32'b10000000000000000111111111110110; // input=-0.84130859375, output=-0.999699514384
			11'd1886: out = 32'b10000000000000001000000000110001; // input=-0.84228515625, output=-1.00150865423
			11'd1887: out = 32'b10000000000000001000000001101101; // input=-0.84326171875, output=-1.00332292294
			11'd1888: out = 32'b10000000000000001000000010101001; // input=-0.84423828125, output=-1.00514237039
			11'd1889: out = 32'b10000000000000001000000011100100; // input=-0.84521484375, output=-1.00696704727
			11'd1890: out = 32'b10000000000000001000000100100000; // input=-0.84619140625, output=-1.00879700506
			11'd1891: out = 32'b10000000000000001000000101011100; // input=-0.84716796875, output=-1.01063229605
			11'd1892: out = 32'b10000000000000001000000110011001; // input=-0.84814453125, output=-1.01247297339
			11'd1893: out = 32'b10000000000000001000000111010101; // input=-0.84912109375, output=-1.01431909107
			11'd1894: out = 32'b10000000000000001000001000010010; // input=-0.85009765625, output=-1.01617070397
			11'd1895: out = 32'b10000000000000001000001001001111; // input=-0.85107421875, output=-1.01802786786
			11'd1896: out = 32'b10000000000000001000001010001100; // input=-0.85205078125, output=-1.01989063942
			11'd1897: out = 32'b10000000000000001000001011001001; // input=-0.85302734375, output=-1.02175907629
			11'd1898: out = 32'b10000000000000001000001100000110; // input=-0.85400390625, output=-1.02363323705
			11'd1899: out = 32'b10000000000000001000001101000100; // input=-0.85498046875, output=-1.02551318129
			11'd1900: out = 32'b10000000000000001000001110000010; // input=-0.85595703125, output=-1.02739896957
			11'd1901: out = 32'b10000000000000001000001111000000; // input=-0.85693359375, output=-1.02929066351
			11'd1902: out = 32'b10000000000000001000001111111110; // input=-0.85791015625, output=-1.03118832579
			11'd1903: out = 32'b10000000000000001000010000111100; // input=-0.85888671875, output=-1.03309202014
			11'd1904: out = 32'b10000000000000001000010001111011; // input=-0.85986328125, output=-1.03500181142
			11'd1905: out = 32'b10000000000000001000010010111010; // input=-0.86083984375, output=-1.03691776563
			11'd1906: out = 32'b10000000000000001000010011111001; // input=-0.86181640625, output=-1.03883994992
			11'd1907: out = 32'b10000000000000001000010100111000; // input=-0.86279296875, output=-1.04076843263
			11'd1908: out = 32'b10000000000000001000010101110111; // input=-0.86376953125, output=-1.04270328333
			11'd1909: out = 32'b10000000000000001000010110110111; // input=-0.86474609375, output=-1.04464457284
			11'd1910: out = 32'b10000000000000001000010111110111; // input=-0.86572265625, output=-1.04659237326
			11'd1911: out = 32'b10000000000000001000011000110111; // input=-0.86669921875, output=-1.04854675801
			11'd1912: out = 32'b10000000000000001000011001110111; // input=-0.86767578125, output=-1.05050780186
			11'd1913: out = 32'b10000000000000001000011010111000; // input=-0.86865234375, output=-1.05247558096
			11'd1914: out = 32'b10000000000000001000011011111000; // input=-0.86962890625, output=-1.0544501729
			11'd1915: out = 32'b10000000000000001000011100111001; // input=-0.87060546875, output=-1.0564316567
			11'd1916: out = 32'b10000000000000001000011101111010; // input=-0.87158203125, output=-1.0584201129
			11'd1917: out = 32'b10000000000000001000011110111100; // input=-0.87255859375, output=-1.06041562356
			11'd1918: out = 32'b10000000000000001000011111111101; // input=-0.87353515625, output=-1.06241827236
			11'd1919: out = 32'b10000000000000001000100000111111; // input=-0.87451171875, output=-1.06442814454
			11'd1920: out = 32'b10000000000000001000100010000001; // input=-0.87548828125, output=-1.06644532706
			11'd1921: out = 32'b10000000000000001000100011000100; // input=-0.87646484375, output=-1.06846990857
			11'd1922: out = 32'b10000000000000001000100100000110; // input=-0.87744140625, output=-1.07050197947
			11'd1923: out = 32'b10000000000000001000100101001001; // input=-0.87841796875, output=-1.07254163199
			11'd1924: out = 32'b10000000000000001000100110001100; // input=-0.87939453125, output=-1.0745889602
			11'd1925: out = 32'b10000000000000001000100111001111; // input=-0.88037109375, output=-1.07664406011
			11'd1926: out = 32'b10000000000000001000101000010011; // input=-0.88134765625, output=-1.07870702967
			11'd1927: out = 32'b10000000000000001000101001010111; // input=-0.88232421875, output=-1.08077796888
			11'd1928: out = 32'b10000000000000001000101010011011; // input=-0.88330078125, output=-1.08285697979
			11'd1929: out = 32'b10000000000000001000101011011111; // input=-0.88427734375, output=-1.08494416663
			11'd1930: out = 32'b10000000000000001000101100100100; // input=-0.88525390625, output=-1.08703963583
			11'd1931: out = 32'b10000000000000001000101101101001; // input=-0.88623046875, output=-1.08914349607
			11'd1932: out = 32'b10000000000000001000101110101110; // input=-0.88720703125, output=-1.09125585841
			11'd1933: out = 32'b10000000000000001000101111110100; // input=-0.88818359375, output=-1.09337683631
			11'd1934: out = 32'b10000000000000001000110000111010; // input=-0.88916015625, output=-1.0955065457
			11'd1935: out = 32'b10000000000000001000110010000000; // input=-0.89013671875, output=-1.0976451051
			11'd1936: out = 32'b10000000000000001000110011000110; // input=-0.89111328125, output=-1.09979263568
			11'd1937: out = 32'b10000000000000001000110100001101; // input=-0.89208984375, output=-1.10194926132
			11'd1938: out = 32'b10000000000000001000110101010100; // input=-0.89306640625, output=-1.10411510871
			11'd1939: out = 32'b10000000000000001000110110011011; // input=-0.89404296875, output=-1.10629030749
			11'd1940: out = 32'b10000000000000001000110111100011; // input=-0.89501953125, output=-1.10847499025
			11'd1941: out = 32'b10000000000000001000111000101010; // input=-0.89599609375, output=-1.1106692927
			11'd1942: out = 32'b10000000000000001000111001110011; // input=-0.89697265625, output=-1.11287335376
			11'd1943: out = 32'b10000000000000001000111010111011; // input=-0.89794921875, output=-1.11508731565
			11'd1944: out = 32'b10000000000000001000111100000100; // input=-0.89892578125, output=-1.117311324
			11'd1945: out = 32'b10000000000000001000111101001101; // input=-0.89990234375, output=-1.11954552799
			11'd1946: out = 32'b10000000000000001000111110010111; // input=-0.90087890625, output=-1.12179008044
			11'd1947: out = 32'b10000000000000001000111111100001; // input=-0.90185546875, output=-1.12404513797
			11'd1948: out = 32'b10000000000000001001000000101011; // input=-0.90283203125, output=-1.1263108611
			11'd1949: out = 32'b10000000000000001001000001110110; // input=-0.90380859375, output=-1.12858741441
			11'd1950: out = 32'b10000000000000001001000011000001; // input=-0.90478515625, output=-1.13087496667
			11'd1951: out = 32'b10000000000000001001000100001100; // input=-0.90576171875, output=-1.13317369102
			11'd1952: out = 32'b10000000000000001001000101011000; // input=-0.90673828125, output=-1.13548376509
			11'd1953: out = 32'b10000000000000001001000110100100; // input=-0.90771484375, output=-1.13780537118
			11'd1954: out = 32'b10000000000000001001000111110000; // input=-0.90869140625, output=-1.14013869645
			11'd1955: out = 32'b10000000000000001001001000111101; // input=-0.90966796875, output=-1.14248393307
			11'd1956: out = 32'b10000000000000001001001010001010; // input=-0.91064453125, output=-1.14484127846
			11'd1957: out = 32'b10000000000000001001001011011000; // input=-0.91162109375, output=-1.14721093543
			11'd1958: out = 32'b10000000000000001001001100100110; // input=-0.91259765625, output=-1.14959311244
			11'd1959: out = 32'b10000000000000001001001101110100; // input=-0.91357421875, output=-1.1519880238
			11'd1960: out = 32'b10000000000000001001001111000011; // input=-0.91455078125, output=-1.1543958899
			11'd1961: out = 32'b10000000000000001001010000010011; // input=-0.91552734375, output=-1.15681693745
			11'd1962: out = 32'b10000000000000001001010001100010; // input=-0.91650390625, output=-1.15925139978
			11'd1963: out = 32'b10000000000000001001010010110011; // input=-0.91748046875, output=-1.16169951703
			11'd1964: out = 32'b10000000000000001001010100000011; // input=-0.91845703125, output=-1.16416153653
			11'd1965: out = 32'b10000000000000001001010101010100; // input=-0.91943359375, output=-1.16663771301
			11'd1966: out = 32'b10000000000000001001010110100110; // input=-0.92041015625, output=-1.16912830899
			11'd1967: out = 32'b10000000000000001001010111111000; // input=-0.92138671875, output=-1.17163359507
			11'd1968: out = 32'b10000000000000001001011001001011; // input=-0.92236328125, output=-1.17415385031
			11'd1969: out = 32'b10000000000000001001011010011110; // input=-0.92333984375, output=-1.17668936258
			11'd1970: out = 32'b10000000000000001001011011110001; // input=-0.92431640625, output=-1.17924042897
			11'd1971: out = 32'b10000000000000001001011101000101; // input=-0.92529296875, output=-1.18180735621
			11'd1972: out = 32'b10000000000000001001011110011010; // input=-0.92626953125, output=-1.1843904611
			11'd1973: out = 32'b10000000000000001001011111101111; // input=-0.92724609375, output=-1.18699007099
			11'd1974: out = 32'b10000000000000001001100001000101; // input=-0.92822265625, output=-1.18960652428
			11'd1975: out = 32'b10000000000000001001100010011011; // input=-0.92919921875, output=-1.19224017094
			11'd1976: out = 32'b10000000000000001001100011110010; // input=-0.93017578125, output=-1.19489137306
			11'd1977: out = 32'b10000000000000001001100101001010; // input=-0.93115234375, output=-1.1975605055
			11'd1978: out = 32'b10000000000000001001100110100010; // input=-0.93212890625, output=-1.20024795643
			11'd1979: out = 32'b10000000000000001001100111111010; // input=-0.93310546875, output=-1.20295412811
			11'd1980: out = 32'b10000000000000001001101001010100; // input=-0.93408203125, output=-1.20567943755
			11'd1981: out = 32'b10000000000000001001101010101110; // input=-0.93505859375, output=-1.20842431728
			11'd1982: out = 32'b10000000000000001001101100001000; // input=-0.93603515625, output=-1.21118921619
			11'd1983: out = 32'b10000000000000001001101101100100; // input=-0.93701171875, output=-1.2139746004
			11'd1984: out = 32'b10000000000000001001101110111111; // input=-0.93798828125, output=-1.21678095422
			11'd1985: out = 32'b10000000000000001001110000011100; // input=-0.93896484375, output=-1.21960878111
			11'd1986: out = 32'b10000000000000001001110001111010; // input=-0.93994140625, output=-1.22245860481
			11'd1987: out = 32'b10000000000000001001110011011000; // input=-0.94091796875, output=-1.22533097047
			11'd1988: out = 32'b10000000000000001001110100110111; // input=-0.94189453125, output=-1.22822644589
			11'd1989: out = 32'b10000000000000001001110110010110; // input=-0.94287109375, output=-1.23114562288
			11'd1990: out = 32'b10000000000000001001110111110111; // input=-0.94384765625, output=-1.23408911871
			11'd1991: out = 32'b10000000000000001001111001011000; // input=-0.94482421875, output=-1.23705757763
			11'd1992: out = 32'b10000000000000001001111010111010; // input=-0.94580078125, output=-1.24005167258
			11'd1993: out = 32'b10000000000000001001111100011101; // input=-0.94677734375, output=-1.24307210702
			11'd1994: out = 32'b10000000000000001001111110000001; // input=-0.94775390625, output=-1.24611961686
			11'd1995: out = 32'b10000000000000001001111111100110; // input=-0.94873046875, output=-1.24919497264
			11'd1996: out = 32'b10000000000000001010000001001011; // input=-0.94970703125, output=-1.25229898181
			11'd1997: out = 32'b10000000000000001010000010110010; // input=-0.95068359375, output=-1.25543249128
			11'd1998: out = 32'b10000000000000001010000100011010; // input=-0.95166015625, output=-1.25859639018
			11'd1999: out = 32'b10000000000000001010000110000010; // input=-0.95263671875, output=-1.26179161284
			11'd2000: out = 32'b10000000000000001010000111101100; // input=-0.95361328125, output=-1.26501914206
			11'd2001: out = 32'b10000000000000001010001001010111; // input=-0.95458984375, output=-1.26828001276
			11'd2002: out = 32'b10000000000000001010001011000011; // input=-0.95556640625, output=-1.27157531586
			11'd2003: out = 32'b10000000000000001010001100110000; // input=-0.95654296875, output=-1.27490620266
			11'd2004: out = 32'b10000000000000001010001110011110; // input=-0.95751953125, output=-1.27827388961
			11'd2005: out = 32'b10000000000000001010010000001110; // input=-0.95849609375, output=-1.28167966359
			11'd2006: out = 32'b10000000000000001010010001111111; // input=-0.95947265625, output=-1.28512488772
			11'd2007: out = 32'b10000000000000001010010011110001; // input=-0.96044921875, output=-1.28861100788
			11'd2008: out = 32'b10000000000000001010010101100101; // input=-0.96142578125, output=-1.2921395599
			11'd2009: out = 32'b10000000000000001010010111011010; // input=-0.96240234375, output=-1.29571217755
			11'd2010: out = 32'b10000000000000001010011001010000; // input=-0.96337890625, output=-1.29933060156
			11'd2011: out = 32'b10000000000000001010011011001001; // input=-0.96435546875, output=-1.30299668967
			11'd2012: out = 32'b10000000000000001010011101000010; // input=-0.96533203125, output=-1.30671242792
			11'd2013: out = 32'b10000000000000001010011110111110; // input=-0.96630859375, output=-1.3104799434
			11'd2014: out = 32'b10000000000000001010100000111011; // input=-0.96728515625, output=-1.31430151869
			11'd2015: out = 32'b10000000000000001010100010111010; // input=-0.96826171875, output=-1.31817960826
			11'd2016: out = 32'b10000000000000001010100100111011; // input=-0.96923828125, output=-1.32211685711
			11'd2017: out = 32'b10000000000000001010100110111110; // input=-0.97021484375, output=-1.32611612215
			11'd2018: out = 32'b10000000000000001010101001000011; // input=-0.97119140625, output=-1.33018049673
			11'd2019: out = 32'b10000000000000001010101011001011; // input=-0.97216796875, output=-1.33431333899
			11'd2020: out = 32'b10000000000000001010101101010101; // input=-0.97314453125, output=-1.33851830468
			11'd2021: out = 32'b10000000000000001010101111100001; // input=-0.97412109375, output=-1.34279938541
			11'd2022: out = 32'b10000000000000001010110001110000; // input=-0.97509765625, output=-1.34716095354
			11'd2023: out = 32'b10000000000000001010110100000001; // input=-0.97607421875, output=-1.35160781497
			11'd2024: out = 32'b10000000000000001010110110010110; // input=-0.97705078125, output=-1.35614527182
			11'd2025: out = 32'b10000000000000001010111000101110; // input=-0.97802734375, output=-1.36077919721
			11'd2026: out = 32'b10000000000000001010111011001001; // input=-0.97900390625, output=-1.36551612523
			11'd2027: out = 32'b10000000000000001010111101101000; // input=-0.97998046875, output=-1.37036335996
			11'd2028: out = 32'b10000000000000001011000000001011; // input=-0.98095703125, output=-1.37532910873
			11'd2029: out = 32'b10000000000000001011000010110010; // input=-0.98193359375, output=-1.38042264672
			11'd2030: out = 32'b10000000000000001011000101011101; // input=-0.98291015625, output=-1.38565452202
			11'd2031: out = 32'b10000000000000001011001000001101; // input=-0.98388671875, output=-1.39103681451
			11'd2032: out = 32'b10000000000000001011001011000011; // input=-0.98486328125, output=-1.39658346647
			11'd2033: out = 32'b10000000000000001011001101111111; // input=-0.98583984375, output=-1.40231071107
			11'd2034: out = 32'b10000000000000001011010001000001; // input=-0.98681640625, output=-1.40823763659
			11'd2035: out = 32'b10000000000000001011010100001011; // input=-0.98779296875, output=-1.41438694293
			11'd2036: out = 32'b10000000000000001011010111011100; // input=-0.98876953125, output=-1.42078597714
			11'd2037: out = 32'b10000000000000001011011010110111; // input=-0.98974609375, output=-1.42746818517
			11'd2038: out = 32'b10000000000000001011011110011101; // input=-0.99072265625, output=-1.43447520447
			11'd2039: out = 32'b10000000000000001011100010001111; // input=-0.99169921875, output=-1.44185998152
			11'd2040: out = 32'b10000000000000001011100110001111; // input=-0.99267578125, output=-1.44969160393
			11'd2041: out = 32'b10000000000000001011101010100010; // input=-0.99365234375, output=-1.45806316311
			11'd2042: out = 32'b10000000000000001011101111001010; // input=-0.99462890625, output=-1.46710535557
			11'd2043: out = 32'b10000000000000001011110100001111; // input=-0.99560546875, output=-1.47701196053
			11'd2044: out = 32'b10000000000000001011111001111010; // input=-0.99658203125, output=-1.48809303047
			11'd2045: out = 32'b10000000000000001100000000011110; // input=-0.99755859375, output=-1.50090497815
			11'd2046: out = 32'b10000000000000001100001000100010; // input=-0.99853515625, output=-1.51666312963
			11'd2047: out = 32'b10000000000000001100010100010000; // input=-0.99951171875, output=-1.53954505509
		endcase
	end
	converter U0 (a, index);

endmodule

module cos_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000000111111111111111; // input=0.001953125, output=0.999998092652
			11'd1: out = 32'b00000000000000000111111111111111; // input=0.005859375, output=0.999982833911
			11'd2: out = 32'b00000000000000000111111111111110; // input=0.009765625, output=0.999952316663
			11'd3: out = 32'b00000000000000000111111111111101; // input=0.013671875, output=0.999906541373
			11'd4: out = 32'b00000000000000000111111111111011; // input=0.017578125, output=0.999845508739
			11'd5: out = 32'b00000000000000000111111111111000; // input=0.021484375, output=0.999769219693
			11'd6: out = 32'b00000000000000000111111111110101; // input=0.025390625, output=0.999677675398
			11'd7: out = 32'b00000000000000000111111111110010; // input=0.029296875, output=0.999570877252
			11'd8: out = 32'b00000000000000000111111111101110; // input=0.033203125, output=0.999448826885
			11'd9: out = 32'b00000000000000000111111111101001; // input=0.037109375, output=0.999311526157
			11'd10: out = 32'b00000000000000000111111111100100; // input=0.041015625, output=0.999158977166
			11'd11: out = 32'b00000000000000000111111111011111; // input=0.044921875, output=0.998991182238
			11'd12: out = 32'b00000000000000000111111111011001; // input=0.048828125, output=0.998808143933
			11'd13: out = 32'b00000000000000000111111111010010; // input=0.052734375, output=0.998609865045
			11'd14: out = 32'b00000000000000000111111111001011; // input=0.056640625, output=0.998396348599
			11'd15: out = 32'b00000000000000000111111111000100; // input=0.060546875, output=0.998167597854
			11'd16: out = 32'b00000000000000000111111110111100; // input=0.064453125, output=0.997923616299
			11'd17: out = 32'b00000000000000000111111110110011; // input=0.068359375, output=0.997664407657
			11'd18: out = 32'b00000000000000000111111110101010; // input=0.072265625, output=0.997389975884
			11'd19: out = 32'b00000000000000000111111110100001; // input=0.076171875, output=0.997100325166
			11'd20: out = 32'b00000000000000000111111110010111; // input=0.080078125, output=0.996795459925
			11'd21: out = 32'b00000000000000000111111110001101; // input=0.083984375, output=0.996475384812
			11'd22: out = 32'b00000000000000000111111110000010; // input=0.087890625, output=0.99614010471
			11'd23: out = 32'b00000000000000000111111101110110; // input=0.091796875, output=0.995789624735
			11'd24: out = 32'b00000000000000000111111101101010; // input=0.095703125, output=0.995423950236
			11'd25: out = 32'b00000000000000000111111101011110; // input=0.099609375, output=0.995043086793
			11'd26: out = 32'b00000000000000000111111101010001; // input=0.103515625, output=0.994647040216
			11'd27: out = 32'b00000000000000000111111101000011; // input=0.107421875, output=0.994235816549
			11'd28: out = 32'b00000000000000000111111100110101; // input=0.111328125, output=0.993809422066
			11'd29: out = 32'b00000000000000000111111100100111; // input=0.115234375, output=0.993367863275
			11'd30: out = 32'b00000000000000000111111100011000; // input=0.119140625, output=0.992911146912
			11'd31: out = 32'b00000000000000000111111100001000; // input=0.123046875, output=0.992439279947
			11'd32: out = 32'b00000000000000000111111011111000; // input=0.126953125, output=0.991952269579
			11'd33: out = 32'b00000000000000000111111011101000; // input=0.130859375, output=0.99145012324
			11'd34: out = 32'b00000000000000000111111011010111; // input=0.134765625, output=0.990932848592
			11'd35: out = 32'b00000000000000000111111011000101; // input=0.138671875, output=0.990400453528
			11'd36: out = 32'b00000000000000000111111010110100; // input=0.142578125, output=0.989852946172
			11'd37: out = 32'b00000000000000000111111010100001; // input=0.146484375, output=0.989290334878
			11'd38: out = 32'b00000000000000000111111010001110; // input=0.150390625, output=0.98871262823
			11'd39: out = 32'b00000000000000000111111001111011; // input=0.154296875, output=0.988119835044
			11'd40: out = 32'b00000000000000000111111001100111; // input=0.158203125, output=0.987511964365
			11'd41: out = 32'b00000000000000000111111001010010; // input=0.162109375, output=0.986889025468
			11'd42: out = 32'b00000000000000000111111000111101; // input=0.166015625, output=0.986251027859
			11'd43: out = 32'b00000000000000000111111000101000; // input=0.169921875, output=0.985597981273
			11'd44: out = 32'b00000000000000000111111000010010; // input=0.173828125, output=0.984929895674
			11'd45: out = 32'b00000000000000000111110111111100; // input=0.177734375, output=0.984246781257
			11'd46: out = 32'b00000000000000000111110111100101; // input=0.181640625, output=0.983548648445
			11'd47: out = 32'b00000000000000000111110111001110; // input=0.185546875, output=0.98283550789
			11'd48: out = 32'b00000000000000000111110110110110; // input=0.189453125, output=0.982107370475
			11'd49: out = 32'b00000000000000000111110110011101; // input=0.193359375, output=0.98136424731
			11'd50: out = 32'b00000000000000000111110110000101; // input=0.197265625, output=0.980606149734
			11'd51: out = 32'b00000000000000000111110101101011; // input=0.201171875, output=0.979833089314
			11'd52: out = 32'b00000000000000000111110101010001; // input=0.205078125, output=0.979045077847
			11'd53: out = 32'b00000000000000000111110100110111; // input=0.208984375, output=0.978242127357
			11'd54: out = 32'b00000000000000000111110100011100; // input=0.212890625, output=0.977424250095
			11'd55: out = 32'b00000000000000000111110100000001; // input=0.216796875, output=0.976591458542
			11'd56: out = 32'b00000000000000000111110011100101; // input=0.220703125, output=0.975743765405
			11'd57: out = 32'b00000000000000000111110011001001; // input=0.224609375, output=0.974881183619
			11'd58: out = 32'b00000000000000000111110010101100; // input=0.228515625, output=0.974003726345
			11'd59: out = 32'b00000000000000000111110010001111; // input=0.232421875, output=0.973111406972
			11'd60: out = 32'b00000000000000000111110001110001; // input=0.236328125, output=0.972204239117
			11'd61: out = 32'b00000000000000000111110001010011; // input=0.240234375, output=0.971282236621
			11'd62: out = 32'b00000000000000000111110000110100; // input=0.244140625, output=0.970345413553
			11'd63: out = 32'b00000000000000000111110000010101; // input=0.248046875, output=0.969393784208
			11'd64: out = 32'b00000000000000000111101111110101; // input=0.251953125, output=0.968427363107
			11'd65: out = 32'b00000000000000000111101111010101; // input=0.255859375, output=0.967446164995
			11'd66: out = 32'b00000000000000000111101110110101; // input=0.259765625, output=0.966450204846
			11'd67: out = 32'b00000000000000000111101110010100; // input=0.263671875, output=0.965439497855
			11'd68: out = 32'b00000000000000000111101101110010; // input=0.267578125, output=0.964414059445
			11'd69: out = 32'b00000000000000000111101101010000; // input=0.271484375, output=0.963373905264
			11'd70: out = 32'b00000000000000000111101100101101; // input=0.275390625, output=0.962319051181
			11'd71: out = 32'b00000000000000000111101100001010; // input=0.279296875, output=0.961249513295
			11'd72: out = 32'b00000000000000000111101011100111; // input=0.283203125, output=0.960165307923
			11'd73: out = 32'b00000000000000000111101011000011; // input=0.287109375, output=0.95906645161
			11'd74: out = 32'b00000000000000000111101010011110; // input=0.291015625, output=0.957952961123
			11'd75: out = 32'b00000000000000000111101001111001; // input=0.294921875, output=0.956824853452
			11'd76: out = 32'b00000000000000000111101001010100; // input=0.298828125, output=0.955682145811
			11'd77: out = 32'b00000000000000000111101000101110; // input=0.302734375, output=0.954524855637
			11'd78: out = 32'b00000000000000000111101000000111; // input=0.306640625, output=0.953353000587
			11'd79: out = 32'b00000000000000000111100111100001; // input=0.310546875, output=0.952166598544
			11'd80: out = 32'b00000000000000000111100110111001; // input=0.314453125, output=0.95096566761
			11'd81: out = 32'b00000000000000000111100110010001; // input=0.318359375, output=0.94975022611
			11'd82: out = 32'b00000000000000000111100101101001; // input=0.322265625, output=0.94852029259
			11'd83: out = 32'b00000000000000000111100101000000; // input=0.326171875, output=0.947275885817
			11'd84: out = 32'b00000000000000000111100100010111; // input=0.330078125, output=0.94601702478
			11'd85: out = 32'b00000000000000000111100011101101; // input=0.333984375, output=0.944743728687
			11'd86: out = 32'b00000000000000000111100011000011; // input=0.337890625, output=0.943456016966
			11'd87: out = 32'b00000000000000000111100010011000; // input=0.341796875, output=0.942153909268
			11'd88: out = 32'b00000000000000000111100001101101; // input=0.345703125, output=0.940837425461
			11'd89: out = 32'b00000000000000000111100001000010; // input=0.349609375, output=0.939506585632
			11'd90: out = 32'b00000000000000000111100000010110; // input=0.353515625, output=0.938161410088
			11'd91: out = 32'b00000000000000000111011111101001; // input=0.357421875, output=0.936801919355
			11'd92: out = 32'b00000000000000000111011110111100; // input=0.361328125, output=0.935428134178
			11'd93: out = 32'b00000000000000000111011110001111; // input=0.365234375, output=0.934040075518
			11'd94: out = 32'b00000000000000000111011101100001; // input=0.369140625, output=0.932637764556
			11'd95: out = 32'b00000000000000000111011100110010; // input=0.373046875, output=0.931221222689
			11'd96: out = 32'b00000000000000000111011100000011; // input=0.376953125, output=0.929790471532
			11'd97: out = 32'b00000000000000000111011011010100; // input=0.380859375, output=0.928345532916
			11'd98: out = 32'b00000000000000000111011010100100; // input=0.384765625, output=0.92688642889
			11'd99: out = 32'b00000000000000000111011001110100; // input=0.388671875, output=0.925413181717
			11'd100: out = 32'b00000000000000000111011001000011; // input=0.392578125, output=0.923925813877
			11'd101: out = 32'b00000000000000000111011000010010; // input=0.396484375, output=0.922424348067
			11'd102: out = 32'b00000000000000000111010111100000; // input=0.400390625, output=0.920908807195
			11'd103: out = 32'b00000000000000000111010110101110; // input=0.404296875, output=0.919379214389
			11'd104: out = 32'b00000000000000000111010101111100; // input=0.408203125, output=0.917835592986
			11'd105: out = 32'b00000000000000000111010101001001; // input=0.412109375, output=0.916277966542
			11'd106: out = 32'b00000000000000000111010100010101; // input=0.416015625, output=0.914706358823
			11'd107: out = 32'b00000000000000000111010011100001; // input=0.419921875, output=0.913120793811
			11'd108: out = 32'b00000000000000000111010010101101; // input=0.423828125, output=0.911521295699
			11'd109: out = 32'b00000000000000000111010001111000; // input=0.427734375, output=0.909907888893
			11'd110: out = 32'b00000000000000000111010001000011; // input=0.431640625, output=0.908280598013
			11'd111: out = 32'b00000000000000000111010000001101; // input=0.435546875, output=0.906639447888
			11'd112: out = 32'b00000000000000000111001111010111; // input=0.439453125, output=0.90498446356
			11'd113: out = 32'b00000000000000000111001110100000; // input=0.443359375, output=0.903315670283
			11'd114: out = 32'b00000000000000000111001101101001; // input=0.447265625, output=0.901633093521
			11'd115: out = 32'b00000000000000000111001100110001; // input=0.451171875, output=0.899936758946
			11'd116: out = 32'b00000000000000000111001011111001; // input=0.455078125, output=0.898226692444
			11'd117: out = 32'b00000000000000000111001011000001; // input=0.458984375, output=0.896502920108
			11'd118: out = 32'b00000000000000000111001010001000; // input=0.462890625, output=0.89476546824
			11'd119: out = 32'b00000000000000000111001001001110; // input=0.466796875, output=0.893014363352
			11'd120: out = 32'b00000000000000000111001000010100; // input=0.470703125, output=0.891249632163
			11'd121: out = 32'b00000000000000000111000111011010; // input=0.474609375, output=0.889471301602
			11'd122: out = 32'b00000000000000000111000110011111; // input=0.478515625, output=0.887679398803
			11'd123: out = 32'b00000000000000000111000101100100; // input=0.482421875, output=0.885873951108
			11'd124: out = 32'b00000000000000000111000100101001; // input=0.486328125, output=0.884054986067
			11'd125: out = 32'b00000000000000000111000011101101; // input=0.490234375, output=0.882222531435
			11'd126: out = 32'b00000000000000000111000010110000; // input=0.494140625, output=0.880376615172
			11'd127: out = 32'b00000000000000000111000001110011; // input=0.498046875, output=0.878517265445
			11'd128: out = 32'b00000000000000000111000000110110; // input=0.501953125, output=0.876644510625
			11'd129: out = 32'b00000000000000000110111111111000; // input=0.505859375, output=0.874758379289
			11'd130: out = 32'b00000000000000000110111110111010; // input=0.509765625, output=0.872858900216
			11'd131: out = 32'b00000000000000000110111101111011; // input=0.513671875, output=0.870946102391
			11'd132: out = 32'b00000000000000000110111100111100; // input=0.517578125, output=0.869020014999
			11'd133: out = 32'b00000000000000000110111011111100; // input=0.521484375, output=0.867080667431
			11'd134: out = 32'b00000000000000000110111010111101; // input=0.525390625, output=0.865128089279
			11'd135: out = 32'b00000000000000000110111001111100; // input=0.529296875, output=0.863162310337
			11'd136: out = 32'b00000000000000000110111000111011; // input=0.533203125, output=0.861183360599
			11'd137: out = 32'b00000000000000000110110111111010; // input=0.537109375, output=0.859191270264
			11'd138: out = 32'b00000000000000000110110110111000; // input=0.541015625, output=0.857186069726
			11'd139: out = 32'b00000000000000000110110101110110; // input=0.544921875, output=0.855167789584
			11'd140: out = 32'b00000000000000000110110100110100; // input=0.548828125, output=0.853136460634
			11'd141: out = 32'b00000000000000000110110011110001; // input=0.552734375, output=0.85109211387
			11'd142: out = 32'b00000000000000000110110010101101; // input=0.556640625, output=0.849034780489
			11'd143: out = 32'b00000000000000000110110001101001; // input=0.560546875, output=0.846964491881
			11'd144: out = 32'b00000000000000000110110000100101; // input=0.564453125, output=0.844881279637
			11'd145: out = 32'b00000000000000000110101111100000; // input=0.568359375, output=0.842785175544
			11'd146: out = 32'b00000000000000000110101110011011; // input=0.572265625, output=0.840676211586
			11'd147: out = 32'b00000000000000000110101101010110; // input=0.576171875, output=0.838554419944
			11'd148: out = 32'b00000000000000000110101100010000; // input=0.580078125, output=0.836419832992
			11'd149: out = 32'b00000000000000000110101011001001; // input=0.583984375, output=0.834272483304
			11'd150: out = 32'b00000000000000000110101010000011; // input=0.587890625, output=0.832112403643
			11'd151: out = 32'b00000000000000000110101000111011; // input=0.591796875, output=0.829939626972
			11'd152: out = 32'b00000000000000000110100111110100; // input=0.595703125, output=0.827754186442
			11'd153: out = 32'b00000000000000000110100110101100; // input=0.599609375, output=0.825556115402
			11'd154: out = 32'b00000000000000000110100101100011; // input=0.603515625, output=0.823345447392
			11'd155: out = 32'b00000000000000000110100100011011; // input=0.607421875, output=0.821122216143
			11'd156: out = 32'b00000000000000000110100011010001; // input=0.611328125, output=0.818886455579
			11'd157: out = 32'b00000000000000000110100010001000; // input=0.615234375, output=0.816638199815
			11'd158: out = 32'b00000000000000000110100000111110; // input=0.619140625, output=0.814377483157
			11'd159: out = 32'b00000000000000000110011111110011; // input=0.623046875, output=0.812104340101
			11'd160: out = 32'b00000000000000000110011110101000; // input=0.626953125, output=0.809818805332
			11'd161: out = 32'b00000000000000000110011101011101; // input=0.630859375, output=0.807520913724
			11'd162: out = 32'b00000000000000000110011100010001; // input=0.634765625, output=0.80521070034
			11'd163: out = 32'b00000000000000000110011011000101; // input=0.638671875, output=0.802888200432
			11'd164: out = 32'b00000000000000000110011001111001; // input=0.642578125, output=0.800553449438
			11'd165: out = 32'b00000000000000000110011000101100; // input=0.646484375, output=0.798206482983
			11'd166: out = 32'b00000000000000000110010111011110; // input=0.650390625, output=0.795847336879
			11'd167: out = 32'b00000000000000000110010110010001; // input=0.654296875, output=0.793476047124
			11'd168: out = 32'b00000000000000000110010101000011; // input=0.658203125, output=0.791092649901
			11'd169: out = 32'b00000000000000000110010011110100; // input=0.662109375, output=0.788697181577
			11'd170: out = 32'b00000000000000000110010010100101; // input=0.666015625, output=0.786289678704
			11'd171: out = 32'b00000000000000000110010001010110; // input=0.669921875, output=0.783870178019
			11'd172: out = 32'b00000000000000000110010000000110; // input=0.673828125, output=0.781438716439
			11'd173: out = 32'b00000000000000000110001110110110; // input=0.677734375, output=0.778995331066
			11'd174: out = 32'b00000000000000000110001101100110; // input=0.681640625, output=0.776540059182
			11'd175: out = 32'b00000000000000000110001100010101; // input=0.685546875, output=0.774072938252
			11'd176: out = 32'b00000000000000000110001011000100; // input=0.689453125, output=0.771594005922
			11'd177: out = 32'b00000000000000000110001001110010; // input=0.693359375, output=0.769103300017
			11'd178: out = 32'b00000000000000000110001000100000; // input=0.697265625, output=0.766600858541
			11'd179: out = 32'b00000000000000000110000111001110; // input=0.701171875, output=0.76408671968
			11'd180: out = 32'b00000000000000000110000101111011; // input=0.705078125, output=0.761560921795
			11'd181: out = 32'b00000000000000000110000100101000; // input=0.708984375, output=0.759023503428
			11'd182: out = 32'b00000000000000000110000011010100; // input=0.712890625, output=0.756474503295
			11'd183: out = 32'b00000000000000000110000010000000; // input=0.716796875, output=0.753913960293
			11'd184: out = 32'b00000000000000000110000000101100; // input=0.720703125, output=0.751341913491
			11'd185: out = 32'b00000000000000000101111111010111; // input=0.724609375, output=0.748758402136
			11'd186: out = 32'b00000000000000000101111110000010; // input=0.728515625, output=0.746163465649
			11'd187: out = 32'b00000000000000000101111100101101; // input=0.732421875, output=0.743557143625
			11'd188: out = 32'b00000000000000000101111011010111; // input=0.736328125, output=0.740939475835
			11'd189: out = 32'b00000000000000000101111010000001; // input=0.740234375, output=0.738310502219
			11'd190: out = 32'b00000000000000000101111000101010; // input=0.744140625, output=0.735670262894
			11'd191: out = 32'b00000000000000000101110111010100; // input=0.748046875, output=0.733018798145
			11'd192: out = 32'b00000000000000000101110101111100; // input=0.751953125, output=0.730356148432
			11'd193: out = 32'b00000000000000000101110100100101; // input=0.755859375, output=0.727682354382
			11'd194: out = 32'b00000000000000000101110011001101; // input=0.759765625, output=0.724997456795
			11'd195: out = 32'b00000000000000000101110001110100; // input=0.763671875, output=0.722301496639
			11'd196: out = 32'b00000000000000000101110000011100; // input=0.767578125, output=0.71959451505
			11'd197: out = 32'b00000000000000000101101111000011; // input=0.771484375, output=0.716876553335
			11'd198: out = 32'b00000000000000000101101101101001; // input=0.775390625, output=0.714147652965
			11'd199: out = 32'b00000000000000000101101100001111; // input=0.779296875, output=0.711407855581
			11'd200: out = 32'b00000000000000000101101010110101; // input=0.783203125, output=0.708657202988
			11'd201: out = 32'b00000000000000000101101001011011; // input=0.787109375, output=0.705895737158
			11'd202: out = 32'b00000000000000000101101000000000; // input=0.791015625, output=0.703123500228
			11'd203: out = 32'b00000000000000000101100110100101; // input=0.794921875, output=0.700340534498
			11'd204: out = 32'b00000000000000000101100101001001; // input=0.798828125, output=0.697546882433
			11'd205: out = 32'b00000000000000000101100011101101; // input=0.802734375, output=0.694742586661
			11'd206: out = 32'b00000000000000000101100010010001; // input=0.806640625, output=0.691927689972
			11'd207: out = 32'b00000000000000000101100000110101; // input=0.810546875, output=0.689102235318
			11'd208: out = 32'b00000000000000000101011111011000; // input=0.814453125, output=0.686266265812
			11'd209: out = 32'b00000000000000000101011101111010; // input=0.818359375, output=0.683419824726
			11'd210: out = 32'b00000000000000000101011100011101; // input=0.822265625, output=0.680562955495
			11'd211: out = 32'b00000000000000000101011010111111; // input=0.826171875, output=0.677695701711
			11'd212: out = 32'b00000000000000000101011001100000; // input=0.830078125, output=0.674818107123
			11'd213: out = 32'b00000000000000000101011000000010; // input=0.833984375, output=0.671930215642
			11'd214: out = 32'b00000000000000000101010110100011; // input=0.837890625, output=0.669032071333
			11'd215: out = 32'b00000000000000000101010101000100; // input=0.841796875, output=0.666123718417
			11'd216: out = 32'b00000000000000000101010011100100; // input=0.845703125, output=0.663205201273
			11'd217: out = 32'b00000000000000000101010010000100; // input=0.849609375, output=0.660276564433
			11'd218: out = 32'b00000000000000000101010000100100; // input=0.853515625, output=0.657337852585
			11'd219: out = 32'b00000000000000000101001111000011; // input=0.857421875, output=0.654389110571
			11'd220: out = 32'b00000000000000000101001101100010; // input=0.861328125, output=0.651430383384
			11'd221: out = 32'b00000000000000000101001100000001; // input=0.865234375, output=0.64846171617
			11'd222: out = 32'b00000000000000000101001010011111; // input=0.869140625, output=0.645483154229
			11'd223: out = 32'b00000000000000000101001000111101; // input=0.873046875, output=0.642494743009
			11'd224: out = 32'b00000000000000000101000111011011; // input=0.876953125, output=0.63949652811
			11'd225: out = 32'b00000000000000000101000101111000; // input=0.880859375, output=0.63648855528
			11'd226: out = 32'b00000000000000000101000100010110; // input=0.884765625, output=0.633470870418
			11'd227: out = 32'b00000000000000000101000010110010; // input=0.888671875, output=0.63044351957
			11'd228: out = 32'b00000000000000000101000001001111; // input=0.892578125, output=0.62740654893
			11'd229: out = 32'b00000000000000000100111111101011; // input=0.896484375, output=0.624360004837
			11'd230: out = 32'b00000000000000000100111110000111; // input=0.900390625, output=0.621303933779
			11'd231: out = 32'b00000000000000000100111100100010; // input=0.904296875, output=0.618238382388
			11'd232: out = 32'b00000000000000000100111010111110; // input=0.908203125, output=0.615163397439
			11'd233: out = 32'b00000000000000000100111001011001; // input=0.912109375, output=0.612079025854
			11'd234: out = 32'b00000000000000000100110111110011; // input=0.916015625, output=0.608985314696
			11'd235: out = 32'b00000000000000000100110110001110; // input=0.919921875, output=0.605882311171
			11'd236: out = 32'b00000000000000000100110100101000; // input=0.923828125, output=0.602770062628
			11'd237: out = 32'b00000000000000000100110011000001; // input=0.927734375, output=0.599648616555
			11'd238: out = 32'b00000000000000000100110001011011; // input=0.931640625, output=0.596518020582
			11'd239: out = 32'b00000000000000000100101111110100; // input=0.935546875, output=0.593378322478
			11'd240: out = 32'b00000000000000000100101110001101; // input=0.939453125, output=0.590229570151
			11'd241: out = 32'b00000000000000000100101100100101; // input=0.943359375, output=0.587071811646
			11'd242: out = 32'b00000000000000000100101010111101; // input=0.947265625, output=0.583905095149
			11'd243: out = 32'b00000000000000000100101001010101; // input=0.951171875, output=0.580729468977
			11'd244: out = 32'b00000000000000000100100111101101; // input=0.955078125, output=0.577544981589
			11'd245: out = 32'b00000000000000000100100110000100; // input=0.958984375, output=0.574351681575
			11'd246: out = 32'b00000000000000000100100100011011; // input=0.962890625, output=0.571149617661
			11'd247: out = 32'b00000000000000000100100010110010; // input=0.966796875, output=0.567938838706
			11'd248: out = 32'b00000000000000000100100001001001; // input=0.970703125, output=0.564719393703
			11'd249: out = 32'b00000000000000000100011111011111; // input=0.974609375, output=0.561491331777
			11'd250: out = 32'b00000000000000000100011101110101; // input=0.978515625, output=0.558254702185
			11'd251: out = 32'b00000000000000000100011100001011; // input=0.982421875, output=0.555009554312
			11'd252: out = 32'b00000000000000000100011010100000; // input=0.986328125, output=0.551755937677
			11'd253: out = 32'b00000000000000000100011000110101; // input=0.990234375, output=0.548493901924
			11'd254: out = 32'b00000000000000000100010111001010; // input=0.994140625, output=0.54522349683
			11'd255: out = 32'b00000000000000000100010101011110; // input=0.998046875, output=0.541944772296
			11'd256: out = 32'b00000000000000000100010011110011; // input=1.001953125, output=0.538657778351
			11'd257: out = 32'b00000000000000000100010010000111; // input=1.005859375, output=0.535362565152
			11'd258: out = 32'b00000000000000000100010000011011; // input=1.009765625, output=0.532059182978
			11'd259: out = 32'b00000000000000000100001110101110; // input=1.013671875, output=0.528747682236
			11'd260: out = 32'b00000000000000000100001101000001; // input=1.017578125, output=0.525428113455
			11'd261: out = 32'b00000000000000000100001011010100; // input=1.021484375, output=0.522100527287
			11'd262: out = 32'b00000000000000000100001001100111; // input=1.025390625, output=0.518764974507
			11'd263: out = 32'b00000000000000000100000111111001; // input=1.029296875, output=0.515421506013
			11'd264: out = 32'b00000000000000000100000110001100; // input=1.033203125, output=0.51207017282
			11'd265: out = 32'b00000000000000000100000100011101; // input=1.037109375, output=0.508711026066
			11'd266: out = 32'b00000000000000000100000010101111; // input=1.041015625, output=0.505344117008
			11'd267: out = 32'b00000000000000000100000001000001; // input=1.044921875, output=0.501969497021
			11'd268: out = 32'b00000000000000000011111111010010; // input=1.048828125, output=0.498587217597
			11'd269: out = 32'b00000000000000000011111101100011; // input=1.052734375, output=0.495197330345
			11'd270: out = 32'b00000000000000000011111011110011; // input=1.056640625, output=0.491799886991
			11'd271: out = 32'b00000000000000000011111010000100; // input=1.060546875, output=0.488394939376
			11'd272: out = 32'b00000000000000000011111000010100; // input=1.064453125, output=0.484982539455
			11'd273: out = 32'b00000000000000000011110110100100; // input=1.068359375, output=0.481562739297
			11'd274: out = 32'b00000000000000000011110100110100; // input=1.072265625, output=0.478135591084
			11'd275: out = 32'b00000000000000000011110011000011; // input=1.076171875, output=0.474701147111
			11'd276: out = 32'b00000000000000000011110001010010; // input=1.080078125, output=0.471259459782
			11'd277: out = 32'b00000000000000000011101111100001; // input=1.083984375, output=0.467810581613
			11'd278: out = 32'b00000000000000000011101101110000; // input=1.087890625, output=0.464354565231
			11'd279: out = 32'b00000000000000000011101011111110; // input=1.091796875, output=0.460891463369
			11'd280: out = 32'b00000000000000000011101010001101; // input=1.095703125, output=0.45742132887
			11'd281: out = 32'b00000000000000000011101000011011; // input=1.099609375, output=0.453944214685
			11'd282: out = 32'b00000000000000000011100110101001; // input=1.103515625, output=0.45046017387
			11'd283: out = 32'b00000000000000000011100100110110; // input=1.107421875, output=0.446969259586
			11'd284: out = 32'b00000000000000000011100011000100; // input=1.111328125, output=0.443471525102
			11'd285: out = 32'b00000000000000000011100001010001; // input=1.115234375, output=0.439967023787
			11'd286: out = 32'b00000000000000000011011111011110; // input=1.119140625, output=0.436455809118
			11'd287: out = 32'b00000000000000000011011101101011; // input=1.123046875, output=0.432937934669
			11'd288: out = 32'b00000000000000000011011011110111; // input=1.126953125, output=0.429413454121
			11'd289: out = 32'b00000000000000000011011010000011; // input=1.130859375, output=0.425882421251
			11'd290: out = 32'b00000000000000000011011000001111; // input=1.134765625, output=0.42234488994
			11'd291: out = 32'b00000000000000000011010110011011; // input=1.138671875, output=0.418800914165
			11'd292: out = 32'b00000000000000000011010100100111; // input=1.142578125, output=0.415250548003
			11'd293: out = 32'b00000000000000000011010010110010; // input=1.146484375, output=0.411693845629
			11'd294: out = 32'b00000000000000000011010000111110; // input=1.150390625, output=0.408130861314
			11'd295: out = 32'b00000000000000000011001111001001; // input=1.154296875, output=0.404561649424
			11'd296: out = 32'b00000000000000000011001101010100; // input=1.158203125, output=0.40098626442
			11'd297: out = 32'b00000000000000000011001011011110; // input=1.162109375, output=0.39740476086
			11'd298: out = 32'b00000000000000000011001001101001; // input=1.166015625, output=0.393817193392
			11'd299: out = 32'b00000000000000000011000111110011; // input=1.169921875, output=0.390223616758
			11'd300: out = 32'b00000000000000000011000101111101; // input=1.173828125, output=0.386624085792
			11'd301: out = 32'b00000000000000000011000100000111; // input=1.177734375, output=0.383018655418
			11'd302: out = 32'b00000000000000000011000010010000; // input=1.181640625, output=0.37940738065
			11'd303: out = 32'b00000000000000000011000000011010; // input=1.185546875, output=0.375790316593
			11'd304: out = 32'b00000000000000000010111110100011; // input=1.189453125, output=0.372167518438
			11'd305: out = 32'b00000000000000000010111100101100; // input=1.193359375, output=0.368539041464
			11'd306: out = 32'b00000000000000000010111010110101; // input=1.197265625, output=0.364904941038
			11'd307: out = 32'b00000000000000000010111000111110; // input=1.201171875, output=0.361265272612
			11'd308: out = 32'b00000000000000000010110111000110; // input=1.205078125, output=0.357620091721
			11'd309: out = 32'b00000000000000000010110101001111; // input=1.208984375, output=0.353969453989
			11'd310: out = 32'b00000000000000000010110011010111; // input=1.212890625, output=0.350313415118
			11'd311: out = 32'b00000000000000000010110001011111; // input=1.216796875, output=0.346652030895
			11'd312: out = 32'b00000000000000000010101111100111; // input=1.220703125, output=0.342985357189
			11'd313: out = 32'b00000000000000000010101101101111; // input=1.224609375, output=0.339313449948
			11'd314: out = 32'b00000000000000000010101011110110; // input=1.228515625, output=0.335636365202
			11'd315: out = 32'b00000000000000000010101001111101; // input=1.232421875, output=0.331954159057
			11'd316: out = 32'b00000000000000000010101000000101; // input=1.236328125, output=0.328266887701
			11'd317: out = 32'b00000000000000000010100110001100; // input=1.240234375, output=0.324574607395
			11'd318: out = 32'b00000000000000000010100100010011; // input=1.244140625, output=0.320877374481
			11'd319: out = 32'b00000000000000000010100010011001; // input=1.248046875, output=0.317175245372
			11'd320: out = 32'b00000000000000000010100000100000; // input=1.251953125, output=0.31346827656
			11'd321: out = 32'b00000000000000000010011110100110; // input=1.255859375, output=0.309756524607
			11'd322: out = 32'b00000000000000000010011100101100; // input=1.259765625, output=0.306040046151
			11'd323: out = 32'b00000000000000000010011010110010; // input=1.263671875, output=0.3023188979
			11'd324: out = 32'b00000000000000000010011000111000; // input=1.267578125, output=0.298593136635
			11'd325: out = 32'b00000000000000000010010110111110; // input=1.271484375, output=0.294862819205
			11'd326: out = 32'b00000000000000000010010101000100; // input=1.275390625, output=0.291128002532
			11'd327: out = 32'b00000000000000000010010011001001; // input=1.279296875, output=0.287388743604
			11'd328: out = 32'b00000000000000000010010001001110; // input=1.283203125, output=0.283645099478
			11'd329: out = 32'b00000000000000000010001111010100; // input=1.287109375, output=0.279897127276
			11'd330: out = 32'b00000000000000000010001101011001; // input=1.291015625, output=0.276144884188
			11'd331: out = 32'b00000000000000000010001011011110; // input=1.294921875, output=0.272388427469
			11'd332: out = 32'b00000000000000000010001001100010; // input=1.298828125, output=0.268627814438
			11'd333: out = 32'b00000000000000000010000111100111; // input=1.302734375, output=0.264863102477
			11'd334: out = 32'b00000000000000000010000101101100; // input=1.306640625, output=0.26109434903
			11'd335: out = 32'b00000000000000000010000011110000; // input=1.310546875, output=0.257321611606
			11'd336: out = 32'b00000000000000000010000001110100; // input=1.314453125, output=0.25354494777
			11'd337: out = 32'b00000000000000000001111111111000; // input=1.318359375, output=0.24976441515
			11'd338: out = 32'b00000000000000000001111101111100; // input=1.322265625, output=0.245980071432
			11'd339: out = 32'b00000000000000000001111100000000; // input=1.326171875, output=0.242191974361
			11'd340: out = 32'b00000000000000000001111010000100; // input=1.330078125, output=0.238400181739
			11'd341: out = 32'b00000000000000000001111000001000; // input=1.333984375, output=0.234604751423
			11'd342: out = 32'b00000000000000000001110110001011; // input=1.337890625, output=0.230805741327
			11'd343: out = 32'b00000000000000000001110100001110; // input=1.341796875, output=0.22700320942
			11'd344: out = 32'b00000000000000000001110010010010; // input=1.345703125, output=0.223197213723
			11'd345: out = 32'b00000000000000000001110000010101; // input=1.349609375, output=0.219387812311
			11'd346: out = 32'b00000000000000000001101110011000; // input=1.353515625, output=0.215575063311
			11'd347: out = 32'b00000000000000000001101100011011; // input=1.357421875, output=0.211759024901
			11'd348: out = 32'b00000000000000000001101010011110; // input=1.361328125, output=0.207939755308
			11'd349: out = 32'b00000000000000000001101000100001; // input=1.365234375, output=0.204117312811
			11'd350: out = 32'b00000000000000000001100110100011; // input=1.369140625, output=0.200291755735
			11'd351: out = 32'b00000000000000000001100100100110; // input=1.373046875, output=0.196463142453
			11'd352: out = 32'b00000000000000000001100010101000; // input=1.376953125, output=0.192631531385
			11'd353: out = 32'b00000000000000000001100000101010; // input=1.380859375, output=0.188796980997
			11'd354: out = 32'b00000000000000000001011110101101; // input=1.384765625, output=0.184959549799
			11'd355: out = 32'b00000000000000000001011100101111; // input=1.388671875, output=0.181119296346
			11'd356: out = 32'b00000000000000000001011010110001; // input=1.392578125, output=0.177276279236
			11'd357: out = 32'b00000000000000000001011000110011; // input=1.396484375, output=0.173430557107
			11'd358: out = 32'b00000000000000000001010110110101; // input=1.400390625, output=0.169582188642
			11'd359: out = 32'b00000000000000000001010100110111; // input=1.404296875, output=0.165731232561
			11'd360: out = 32'b00000000000000000001010010111000; // input=1.408203125, output=0.161877747625
			11'd361: out = 32'b00000000000000000001010000111010; // input=1.412109375, output=0.158021792634
			11'd362: out = 32'b00000000000000000001001110111100; // input=1.416015625, output=0.154163426425
			11'd363: out = 32'b00000000000000000001001100111101; // input=1.419921875, output=0.150302707872
			11'd364: out = 32'b00000000000000000001001010111111; // input=1.423828125, output=0.146439695884
			11'd365: out = 32'b00000000000000000001001001000000; // input=1.427734375, output=0.142574449407
			11'd366: out = 32'b00000000000000000001000111000001; // input=1.431640625, output=0.138707027419
			11'd367: out = 32'b00000000000000000001000101000010; // input=1.435546875, output=0.134837488933
			11'd368: out = 32'b00000000000000000001000011000011; // input=1.439453125, output=0.130965892992
			11'd369: out = 32'b00000000000000000001000001000101; // input=1.443359375, output=0.127092298673
			11'd370: out = 32'b00000000000000000000111111000110; // input=1.447265625, output=0.123216765082
			11'd371: out = 32'b00000000000000000000111101000111; // input=1.451171875, output=0.119339351355
			11'd372: out = 32'b00000000000000000000111011000111; // input=1.455078125, output=0.115460116656
			11'd373: out = 32'b00000000000000000000111001001000; // input=1.458984375, output=0.111579120177
			11'd374: out = 32'b00000000000000000000110111001001; // input=1.462890625, output=0.107696421139
			11'd375: out = 32'b00000000000000000000110101001010; // input=1.466796875, output=0.103812078785
			11'd376: out = 32'b00000000000000000000110011001010; // input=1.470703125, output=0.0999261523872
			11'd377: out = 32'b00000000000000000000110001001011; // input=1.474609375, output=0.0960387012391
			11'd378: out = 32'b00000000000000000000101111001100; // input=1.478515625, output=0.0921497846586
			11'd379: out = 32'b00000000000000000000101101001100; // input=1.482421875, output=0.0882594619857
			11'd380: out = 32'b00000000000000000000101011001101; // input=1.486328125, output=0.084367792582
			11'd381: out = 32'b00000000000000000000101001001101; // input=1.490234375, output=0.0804748358296
			11'd382: out = 32'b00000000000000000000100111001101; // input=1.494140625, output=0.0765806511302
			11'd383: out = 32'b00000000000000000000100101001110; // input=1.498046875, output=0.0726852979043
			11'd384: out = 32'b00000000000000000000100011001110; // input=1.501953125, output=0.0687888355902
			11'd385: out = 32'b00000000000000000000100001001110; // input=1.505859375, output=0.0648913236431
			11'd386: out = 32'b00000000000000000000011111001111; // input=1.509765625, output=0.0609928215342
			11'd387: out = 32'b00000000000000000000011101001111; // input=1.513671875, output=0.0570933887499
			11'd388: out = 32'b00000000000000000000011011001111; // input=1.517578125, output=0.0531930847907
			11'd389: out = 32'b00000000000000000000011001001111; // input=1.521484375, output=0.0492919691706
			11'd390: out = 32'b00000000000000000000010111001111; // input=1.525390625, output=0.0453901014156
			11'd391: out = 32'b00000000000000000000010101001111; // input=1.529296875, output=0.0414875410635
			11'd392: out = 32'b00000000000000000000010011010000; // input=1.533203125, output=0.0375843476626
			11'd393: out = 32'b00000000000000000000010001010000; // input=1.537109375, output=0.0336805807707
			11'd394: out = 32'b00000000000000000000001111010000; // input=1.541015625, output=0.0297762999547
			11'd395: out = 32'b00000000000000000000001101010000; // input=1.544921875, output=0.0258715647889
			11'd396: out = 32'b00000000000000000000001011010000; // input=1.548828125, output=0.0219664348549
			11'd397: out = 32'b00000000000000000000001001010000; // input=1.552734375, output=0.0180609697401
			11'd398: out = 32'b00000000000000000000000111010000; // input=1.556640625, output=0.0141552290372
			11'd399: out = 32'b00000000000000000000000101010000; // input=1.560546875, output=0.0102492723429
			11'd400: out = 32'b00000000000000000000000011010000; // input=1.564453125, output=0.00634315925725
			11'd401: out = 32'b00000000000000000000000001010000; // input=1.568359375, output=0.00243694938283
			11'd402: out = 32'b10000000000000000000000000110000; // input=1.572265625, output=-0.00146929767644
			11'd403: out = 32'b10000000000000000000000010110000; // input=1.576171875, output=-0.00537552231604
			11'd404: out = 32'b10000000000000000000000100110000; // input=1.580078125, output=-0.00928166493177
			11'd405: out = 32'b10000000000000000000000110110000; // input=1.583984375, output=-0.0131876659207
			11'd406: out = 32'b10000000000000000000001000110000; // input=1.587890625, output=-0.0170934656821
			11'd407: out = 32'b10000000000000000000001010110000; // input=1.591796875, output=-0.0209990046183
			11'd408: out = 32'b10000000000000000000001100110000; // input=1.595703125, output=-0.0249042231354
			11'd409: out = 32'b10000000000000000000001110110000; // input=1.599609375, output=-0.0288090616448
			11'd410: out = 32'b10000000000000000000010000110000; // input=1.603515625, output=-0.0327134605633
			11'd411: out = 32'b10000000000000000000010010110000; // input=1.607421875, output=-0.0366173603147
			11'd412: out = 32'b10000000000000000000010100110000; // input=1.611328125, output=-0.0405207013302
			11'd413: out = 32'b10000000000000000000010110110000; // input=1.615234375, output=-0.0444234240496
			11'd414: out = 32'b10000000000000000000011000110000; // input=1.619140625, output=-0.0483254689223
			11'd415: out = 32'b10000000000000000000011010101111; // input=1.623046875, output=-0.0522267764077
			11'd416: out = 32'b10000000000000000000011100101111; // input=1.626953125, output=-0.0561272869768
			11'd417: out = 32'b10000000000000000000011110101111; // input=1.630859375, output=-0.0600269411126
			11'd418: out = 32'b10000000000000000000100000101111; // input=1.634765625, output=-0.0639256793111
			11'd419: out = 32'b10000000000000000000100010101110; // input=1.638671875, output=-0.0678234420824
			11'd420: out = 32'b10000000000000000000100100101110; // input=1.642578125, output=-0.0717201699514
			11'd421: out = 32'b10000000000000000000100110101110; // input=1.646484375, output=-0.0756158034588
			11'd422: out = 32'b10000000000000000000101000101101; // input=1.650390625, output=-0.0795102831621
			11'd423: out = 32'b10000000000000000000101010101101; // input=1.654296875, output=-0.0834035496363
			11'd424: out = 32'b10000000000000000000101100101101; // input=1.658203125, output=-0.087295543475
			11'd425: out = 32'b10000000000000000000101110101100; // input=1.662109375, output=-0.0911862052911
			11'd426: out = 32'b10000000000000000000110000101011; // input=1.666015625, output=-0.0950754757179
			11'd427: out = 32'b10000000000000000000110010101011; // input=1.669921875, output=-0.0989632954099
			11'd428: out = 32'b10000000000000000000110100101010; // input=1.673828125, output=-0.102849605044
			11'd429: out = 32'b10000000000000000000110110101001; // input=1.677734375, output=-0.106734345319
			11'd430: out = 32'b10000000000000000000111000101001; // input=1.681640625, output=-0.11061745696
			11'd431: out = 32'b10000000000000000000111010101000; // input=1.685546875, output=-0.114498880714
			11'd432: out = 32'b10000000000000000000111100100111; // input=1.689453125, output=-0.118378557356
			11'd433: out = 32'b10000000000000000000111110100110; // input=1.693359375, output=-0.122256427688
			11'd434: out = 32'b10000000000000000001000000100101; // input=1.697265625, output=-0.126132432536
			11'd435: out = 32'b10000000000000000001000010100100; // input=1.701171875, output=-0.130006512759
			11'd436: out = 32'b10000000000000000001000100100011; // input=1.705078125, output=-0.133878609242
			11'd437: out = 32'b10000000000000000001000110100010; // input=1.708984375, output=-0.137748662903
			11'd438: out = 32'b10000000000000000001001000100000; // input=1.712890625, output=-0.141616614688
			11'd439: out = 32'b10000000000000000001001010011111; // input=1.716796875, output=-0.145482405578
			11'd440: out = 32'b10000000000000000001001100011110; // input=1.720703125, output=-0.149345976585
			11'd441: out = 32'b10000000000000000001001110011100; // input=1.724609375, output=-0.153207268757
			11'd442: out = 32'b10000000000000000001010000011011; // input=1.728515625, output=-0.157066223174
			11'd443: out = 32'b10000000000000000001010010011001; // input=1.732421875, output=-0.160922780954
			11'd444: out = 32'b10000000000000000001010100010111; // input=1.736328125, output=-0.164776883251
			11'd445: out = 32'b10000000000000000001010110010110; // input=1.740234375, output=-0.168628471254
			11'd446: out = 32'b10000000000000000001011000010100; // input=1.744140625, output=-0.172477486195
			11'd447: out = 32'b10000000000000000001011010010010; // input=1.748046875, output=-0.176323869342
			11'd448: out = 32'b10000000000000000001011100010000; // input=1.751953125, output=-0.180167562003
			11'd449: out = 32'b10000000000000000001011110001110; // input=1.755859375, output=-0.184008505529
			11'd450: out = 32'b10000000000000000001100000001011; // input=1.759765625, output=-0.187846641311
			11'd451: out = 32'b10000000000000000001100010001001; // input=1.763671875, output=-0.191681910785
			11'd452: out = 32'b10000000000000000001100100000111; // input=1.767578125, output=-0.195514255429
			11'd453: out = 32'b10000000000000000001100110000100; // input=1.771484375, output=-0.199343616766
			11'd454: out = 32'b10000000000000000001101000000001; // input=1.775390625, output=-0.203169936364
			11'd455: out = 32'b10000000000000000001101001111111; // input=1.779296875, output=-0.206993155839
			11'd456: out = 32'b10000000000000000001101011111100; // input=1.783203125, output=-0.210813216853
			11'd457: out = 32'b10000000000000000001101101111001; // input=1.787109375, output=-0.214630061117
			11'd458: out = 32'b10000000000000000001101111110110; // input=1.791015625, output=-0.218443630391
			11'd459: out = 32'b10000000000000000001110001110011; // input=1.794921875, output=-0.222253866483
			11'd460: out = 32'b10000000000000000001110011110000; // input=1.798828125, output=-0.226060711255
			11'd461: out = 32'b10000000000000000001110101101100; // input=1.802734375, output=-0.229864106618
			11'd462: out = 32'b10000000000000000001110111101001; // input=1.806640625, output=-0.233663994538
			11'd463: out = 32'b10000000000000000001111001100101; // input=1.810546875, output=-0.237460317033
			11'd464: out = 32'b10000000000000000001111011100001; // input=1.814453125, output=-0.241253016175
			11'd465: out = 32'b10000000000000000001111101011110; // input=1.818359375, output=-0.245042034094
			11'd466: out = 32'b10000000000000000001111111011010; // input=1.822265625, output=-0.248827312972
			11'd467: out = 32'b10000000000000000010000001010101; // input=1.826171875, output=-0.252608795052
			11'd468: out = 32'b10000000000000000010000011010001; // input=1.830078125, output=-0.256386422632
			11'd469: out = 32'b10000000000000000010000101001101; // input=1.833984375, output=-0.260160138071
			11'd470: out = 32'b10000000000000000010000111001000; // input=1.837890625, output=-0.263929883786
			11'd471: out = 32'b10000000000000000010001001000100; // input=1.841796875, output=-0.267695602256
			11'd472: out = 32'b10000000000000000010001010111111; // input=1.845703125, output=-0.271457236021
			11'd473: out = 32'b10000000000000000010001100111010; // input=1.849609375, output=-0.275214727682
			11'd474: out = 32'b10000000000000000010001110110101; // input=1.853515625, output=-0.278968019905
			11'd475: out = 32'b10000000000000000010010000110000; // input=1.857421875, output=-0.282717055419
			11'd476: out = 32'b10000000000000000010010010101011; // input=1.861328125, output=-0.286461777019
			11'd477: out = 32'b10000000000000000010010100100101; // input=1.865234375, output=-0.290202127564
			11'd478: out = 32'b10000000000000000010010110100000; // input=1.869140625, output=-0.293938049982
			11'd479: out = 32'b10000000000000000010011000011010; // input=1.873046875, output=-0.297669487267
			11'd480: out = 32'b10000000000000000010011010010100; // input=1.876953125, output=-0.301396382482
			11'd481: out = 32'b10000000000000000010011100001110; // input=1.880859375, output=-0.305118678759
			11'd482: out = 32'b10000000000000000010011110001000; // input=1.884765625, output=-0.308836319301
			11'd483: out = 32'b10000000000000000010100000000010; // input=1.888671875, output=-0.31254924738
			11'd484: out = 32'b10000000000000000010100001111011; // input=1.892578125, output=-0.316257406342
			11'd485: out = 32'b10000000000000000010100011110100; // input=1.896484375, output=-0.319960739605
			11'd486: out = 32'b10000000000000000010100101101110; // input=1.900390625, output=-0.323659190661
			11'd487: out = 32'b10000000000000000010100111100111; // input=1.904296875, output=-0.327352703076
			11'd488: out = 32'b10000000000000000010101001100000; // input=1.908203125, output=-0.331041220491
			11'd489: out = 32'b10000000000000000010101011011000; // input=1.912109375, output=-0.334724686625
			11'd490: out = 32'b10000000000000000010101101010001; // input=1.916015625, output=-0.338403045272
			11'd491: out = 32'b10000000000000000010101111001001; // input=1.919921875, output=-0.342076240304
			11'd492: out = 32'b10000000000000000010110001000001; // input=1.923828125, output=-0.345744215674
			11'd493: out = 32'b10000000000000000010110010111001; // input=1.927734375, output=-0.349406915413
			11'd494: out = 32'b10000000000000000010110100110001; // input=1.931640625, output=-0.353064283632
			11'd495: out = 32'b10000000000000000010110110101001; // input=1.935546875, output=-0.356716264525
			11'd496: out = 32'b10000000000000000010111000100000; // input=1.939453125, output=-0.360362802366
			11'd497: out = 32'b10000000000000000010111010011000; // input=1.943359375, output=-0.364003841514
			11'd498: out = 32'b10000000000000000010111100001111; // input=1.947265625, output=-0.367639326412
			11'd499: out = 32'b10000000000000000010111110000110; // input=1.951171875, output=-0.371269201585
			11'd500: out = 32'b10000000000000000010111111111101; // input=1.955078125, output=-0.374893411648
			11'd501: out = 32'b10000000000000000011000001110011; // input=1.958984375, output=-0.378511901298
			11'd502: out = 32'b10000000000000000011000011101001; // input=1.962890625, output=-0.382124615322
			11'd503: out = 32'b10000000000000000011000101100000; // input=1.966796875, output=-0.385731498595
			11'd504: out = 32'b10000000000000000011000111010110; // input=1.970703125, output=-0.38933249608
			11'd505: out = 32'b10000000000000000011001001001011; // input=1.974609375, output=-0.392927552829
			11'd506: out = 32'b10000000000000000011001011000001; // input=1.978515625, output=-0.396516613988
			11'd507: out = 32'b10000000000000000011001100110110; // input=1.982421875, output=-0.400099624791
			11'd508: out = 32'b10000000000000000011001110101100; // input=1.986328125, output=-0.403676530566
			11'd509: out = 32'b10000000000000000011010000100001; // input=1.990234375, output=-0.407247276734
			11'd510: out = 32'b10000000000000000011010010010101; // input=1.994140625, output=-0.41081180881
			11'd511: out = 32'b10000000000000000011010100001010; // input=1.998046875, output=-0.414370072403
			11'd512: out = 32'b10000000000000000011010101111110; // input=2.001953125, output=-0.417922013218
			11'd513: out = 32'b10000000000000000011010111110011; // input=2.005859375, output=-0.421467577057
			11'd514: out = 32'b10000000000000000011011001100111; // input=2.009765625, output=-0.42500670982
			11'd515: out = 32'b10000000000000000011011011011010; // input=2.013671875, output=-0.428539357504
			11'd516: out = 32'b10000000000000000011011101001110; // input=2.017578125, output=-0.432065466204
			11'd517: out = 32'b10000000000000000011011111000001; // input=2.021484375, output=-0.435584982116
			11'd518: out = 32'b10000000000000000011100000110100; // input=2.025390625, output=-0.439097851538
			11'd519: out = 32'b10000000000000000011100010100111; // input=2.029296875, output=-0.442604020867
			11'd520: out = 32'b10000000000000000011100100011010; // input=2.033203125, output=-0.446103436603
			11'd521: out = 32'b10000000000000000011100110001100; // input=2.037109375, output=-0.449596045349
			11'd522: out = 32'b10000000000000000011100111111111; // input=2.041015625, output=-0.453081793813
			11'd523: out = 32'b10000000000000000011101001110001; // input=2.044921875, output=-0.456560628806
			11'd524: out = 32'b10000000000000000011101011100010; // input=2.048828125, output=-0.460032497246
			11'd525: out = 32'b10000000000000000011101101010100; // input=2.052734375, output=-0.463497346155
			11'd526: out = 32'b10000000000000000011101111000101; // input=2.056640625, output=-0.466955122666
			11'd527: out = 32'b10000000000000000011110000110110; // input=2.060546875, output=-0.470405774016
			11'd528: out = 32'b10000000000000000011110010100111; // input=2.064453125, output=-0.473849247552
			11'd529: out = 32'b10000000000000000011110100011000; // input=2.068359375, output=-0.477285490732
			11'd530: out = 32'b10000000000000000011110110001000; // input=2.072265625, output=-0.480714451123
			11'd531: out = 32'b10000000000000000011110111111000; // input=2.076171875, output=-0.484136076402
			11'd532: out = 32'b10000000000000000011111001101000; // input=2.080078125, output=-0.487550314361
			11'd533: out = 32'b10000000000000000011111011011000; // input=2.083984375, output=-0.490957112901
			11'd534: out = 32'b10000000000000000011111101000111; // input=2.087890625, output=-0.49435642004
			11'd535: out = 32'b10000000000000000011111110110110; // input=2.091796875, output=-0.497748183909
			11'd536: out = 32'b10000000000000000100000000100101; // input=2.095703125, output=-0.501132352752
			11'd537: out = 32'b10000000000000000100000010010100; // input=2.099609375, output=-0.504508874933
			11'd538: out = 32'b10000000000000000100000100000010; // input=2.103515625, output=-0.507877698929
			11'd539: out = 32'b10000000000000000100000101110000; // input=2.107421875, output=-0.511238773335
			11'd540: out = 32'b10000000000000000100000111011110; // input=2.111328125, output=-0.514592046868
			11'd541: out = 32'b10000000000000000100001001001100; // input=2.115234375, output=-0.517937468358
			11'd542: out = 32'b10000000000000000100001010111001; // input=2.119140625, output=-0.52127498676
			11'd543: out = 32'b10000000000000000100001100100110; // input=2.123046875, output=-0.524604551148
			11'd544: out = 32'b10000000000000000100001110010011; // input=2.126953125, output=-0.527926110715
			11'd545: out = 32'b10000000000000000100010000000000; // input=2.130859375, output=-0.531239614779
			11'd546: out = 32'b10000000000000000100010001101100; // input=2.134765625, output=-0.53454501278
			11'd547: out = 32'b10000000000000000100010011011000; // input=2.138671875, output=-0.537842254283
			11'd548: out = 32'b10000000000000000100010101000100; // input=2.142578125, output=-0.541131288974
			11'd549: out = 32'b10000000000000000100010110101111; // input=2.146484375, output=-0.544412066667
			11'd550: out = 32'b10000000000000000100011000011011; // input=2.150390625, output=-0.547684537302
			11'd551: out = 32'b10000000000000000100011010000101; // input=2.154296875, output=-0.550948650945
			11'd552: out = 32'b10000000000000000100011011110000; // input=2.158203125, output=-0.554204357789
			11'd553: out = 32'b10000000000000000100011101011011; // input=2.162109375, output=-0.557451608157
			11'd554: out = 32'b10000000000000000100011111000101; // input=2.166015625, output=-0.560690352499
			11'd555: out = 32'b10000000000000000100100000101111; // input=2.169921875, output=-0.563920541396
			11'd556: out = 32'b10000000000000000100100010011000; // input=2.173828125, output=-0.567142125559
			11'd557: out = 32'b10000000000000000100100100000001; // input=2.177734375, output=-0.570355055831
			11'd558: out = 32'b10000000000000000100100101101010; // input=2.181640625, output=-0.573559283187
			11'd559: out = 32'b10000000000000000100100111010011; // input=2.185546875, output=-0.576754758734
			11'd560: out = 32'b10000000000000000100101000111100; // input=2.189453125, output=-0.579941433713
			11'd561: out = 32'b10000000000000000100101010100100; // input=2.193359375, output=-0.583119259499
			11'd562: out = 32'b10000000000000000100101100001011; // input=2.197265625, output=-0.586288187603
			11'd563: out = 32'b10000000000000000100101101110011; // input=2.201171875, output=-0.58944816967
			11'd564: out = 32'b10000000000000000100101111011010; // input=2.205078125, output=-0.592599157484
			11'd565: out = 32'b10000000000000000100110001000001; // input=2.208984375, output=-0.595741102963
			11'd566: out = 32'b10000000000000000100110010101000; // input=2.212890625, output=-0.598873958166
			11'd567: out = 32'b10000000000000000100110100001110; // input=2.216796875, output=-0.601997675289
			11'd568: out = 32'b10000000000000000100110101110100; // input=2.220703125, output=-0.605112206669
			11'd569: out = 32'b10000000000000000100110111011010; // input=2.224609375, output=-0.60821750478
			11'd570: out = 32'b10000000000000000100111001000000; // input=2.228515625, output=-0.611313522241
			11'd571: out = 32'b10000000000000000100111010100101; // input=2.232421875, output=-0.61440021181
			11'd572: out = 32'b10000000000000000100111100001010; // input=2.236328125, output=-0.617477526387
			11'd573: out = 32'b10000000000000000100111101101110; // input=2.240234375, output=-0.620545419017
			11'd574: out = 32'b10000000000000000100111111010010; // input=2.244140625, output=-0.623603842888
			11'd575: out = 32'b10000000000000000101000000110110; // input=2.248046875, output=-0.626652751331
			11'd576: out = 32'b10000000000000000101000010011010; // input=2.251953125, output=-0.629692097824
			11'd577: out = 32'b10000000000000000101000011111101; // input=2.255859375, output=-0.63272183599
			11'd578: out = 32'b10000000000000000101000101100000; // input=2.259765625, output=-0.635741919599
			11'd579: out = 32'b10000000000000000101000111000011; // input=2.263671875, output=-0.638752302569
			11'd580: out = 32'b10000000000000000101001000100101; // input=2.267578125, output=-0.641752938965
			11'd581: out = 32'b10000000000000000101001010000111; // input=2.271484375, output=-0.644743783001
			11'd582: out = 32'b10000000000000000101001011101001; // input=2.275390625, output=-0.647724789039
			11'd583: out = 32'b10000000000000000101001101001010; // input=2.279296875, output=-0.650695911595
			11'd584: out = 32'b10000000000000000101001110101011; // input=2.283203125, output=-0.653657105331
			11'd585: out = 32'b10000000000000000101010000001100; // input=2.287109375, output=-0.656608325064
			11'd586: out = 32'b10000000000000000101010001101100; // input=2.291015625, output=-0.659549525762
			11'd587: out = 32'b10000000000000000101010011001100; // input=2.294921875, output=-0.662480662545
			11'd588: out = 32'b10000000000000000101010100101100; // input=2.298828125, output=-0.665401690689
			11'd589: out = 32'b10000000000000000101010110001011; // input=2.302734375, output=-0.668312565622
			11'd590: out = 32'b10000000000000000101010111101010; // input=2.306640625, output=-0.671213242927
			11'd591: out = 32'b10000000000000000101011001001001; // input=2.310546875, output=-0.674103678343
			11'd592: out = 32'b10000000000000000101011010100111; // input=2.314453125, output=-0.676983827767
			11'd593: out = 32'b10000000000000000101011100000101; // input=2.318359375, output=-0.679853647251
			11'd594: out = 32'b10000000000000000101011101100011; // input=2.322265625, output=-0.682713093005
			11'd595: out = 32'b10000000000000000101011111000000; // input=2.326171875, output=-0.685562121397
			11'd596: out = 32'b10000000000000000101100000011110; // input=2.330078125, output=-0.688400688954
			11'd597: out = 32'b10000000000000000101100001111010; // input=2.333984375, output=-0.691228752363
			11'd598: out = 32'b10000000000000000101100011010111; // input=2.337890625, output=-0.694046268473
			11'd599: out = 32'b10000000000000000101100100110010; // input=2.341796875, output=-0.69685319429
			11'd600: out = 32'b10000000000000000101100110001110; // input=2.345703125, output=-0.699649486985
			11'd601: out = 32'b10000000000000000101100111101001; // input=2.349609375, output=-0.702435103889
			11'd602: out = 32'b10000000000000000101101001000100; // input=2.353515625, output=-0.705210002498
			11'd603: out = 32'b10000000000000000101101010011111; // input=2.357421875, output=-0.707974140471
			11'd604: out = 32'b10000000000000000101101011111001; // input=2.361328125, output=-0.710727475628
			11'd605: out = 32'b10000000000000000101101101010011; // input=2.365234375, output=-0.713469965959
			11'd606: out = 32'b10000000000000000101101110101100; // input=2.369140625, output=-0.716201569616
			11'd607: out = 32'b10000000000000000101110000000110; // input=2.373046875, output=-0.718922244918
			11'd608: out = 32'b10000000000000000101110001011110; // input=2.376953125, output=-0.721631950352
			11'd609: out = 32'b10000000000000000101110010110111; // input=2.380859375, output=-0.724330644569
			11'd610: out = 32'b10000000000000000101110100001111; // input=2.384765625, output=-0.727018286392
			11'd611: out = 32'b10000000000000000101110101100111; // input=2.388671875, output=-0.729694834811
			11'd612: out = 32'b10000000000000000101110110111110; // input=2.392578125, output=-0.732360248984
			11'd613: out = 32'b10000000000000000101111000010101; // input=2.396484375, output=-0.735014488241
			11'd614: out = 32'b10000000000000000101111001101100; // input=2.400390625, output=-0.737657512081
			11'd615: out = 32'b10000000000000000101111011000010; // input=2.404296875, output=-0.740289280175
			11'd616: out = 32'b10000000000000000101111100011000; // input=2.408203125, output=-0.742909752365
			11'd617: out = 32'b10000000000000000101111101101101; // input=2.412109375, output=-0.745518888667
			11'd618: out = 32'b10000000000000000101111111000010; // input=2.416015625, output=-0.748116649267
			11'd619: out = 32'b10000000000000000110000000010111; // input=2.419921875, output=-0.750702994528
			11'd620: out = 32'b10000000000000000110000001101011; // input=2.423828125, output=-0.753277884985
			11'd621: out = 32'b10000000000000000110000010111111; // input=2.427734375, output=-0.755841281348
			11'd622: out = 32'b10000000000000000110000100010011; // input=2.431640625, output=-0.758393144503
			11'd623: out = 32'b10000000000000000110000101100110; // input=2.435546875, output=-0.760933435512
			11'd624: out = 32'b10000000000000000110000110111001; // input=2.439453125, output=-0.763462115613
			11'd625: out = 32'b10000000000000000110001000001100; // input=2.443359375, output=-0.765979146221
			11'd626: out = 32'b10000000000000000110001001011110; // input=2.447265625, output=-0.76848448893
			11'd627: out = 32'b10000000000000000110001010101111; // input=2.451171875, output=-0.770978105511
			11'd628: out = 32'b10000000000000000110001100000001; // input=2.455078125, output=-0.773459957915
			11'd629: out = 32'b10000000000000000110001101010010; // input=2.458984375, output=-0.775930008271
			11'd630: out = 32'b10000000000000000110001110100010; // input=2.462890625, output=-0.77838821889
			11'd631: out = 32'b10000000000000000110001111110010; // input=2.466796875, output=-0.780834552263
			11'd632: out = 32'b10000000000000000110010001000010; // input=2.470703125, output=-0.783268971061
			11'd633: out = 32'b10000000000000000110010010010010; // input=2.474609375, output=-0.785691438138
			11'd634: out = 32'b10000000000000000110010011100001; // input=2.478515625, output=-0.78810191653
			11'd635: out = 32'b10000000000000000110010100101111; // input=2.482421875, output=-0.790500369457
			11'd636: out = 32'b10000000000000000110010101111101; // input=2.486328125, output=-0.792886760321
			11'd637: out = 32'b10000000000000000110010111001011; // input=2.490234375, output=-0.795261052708
			11'd638: out = 32'b10000000000000000110011000011001; // input=2.494140625, output=-0.797623210391
			11'd639: out = 32'b10000000000000000110011001100110; // input=2.498046875, output=-0.799973197324
			11'd640: out = 32'b10000000000000000110011010110010; // input=2.501953125, output=-0.802310977651
			11'd641: out = 32'b10000000000000000110011011111110; // input=2.505859375, output=-0.804636515699
			11'd642: out = 32'b10000000000000000110011101001010; // input=2.509765625, output=-0.806949775984
			11'd643: out = 32'b10000000000000000110011110010110; // input=2.513671875, output=-0.809250723208
			11'd644: out = 32'b10000000000000000110011111100001; // input=2.517578125, output=-0.811539322262
			11'd645: out = 32'b10000000000000000110100000101011; // input=2.521484375, output=-0.813815538224
			11'd646: out = 32'b10000000000000000110100001110101; // input=2.525390625, output=-0.816079336362
			11'd647: out = 32'b10000000000000000110100010111111; // input=2.529296875, output=-0.818330682134
			11'd648: out = 32'b10000000000000000110100100001000; // input=2.533203125, output=-0.820569541186
			11'd649: out = 32'b10000000000000000110100101010001; // input=2.537109375, output=-0.822795879357
			11'd650: out = 32'b10000000000000000110100110011010; // input=2.541015625, output=-0.825009662675
			11'd651: out = 32'b10000000000000000110100111100010; // input=2.544921875, output=-0.82721085736
			11'd652: out = 32'b10000000000000000110101000101010; // input=2.548828125, output=-0.829399429826
			11'd653: out = 32'b10000000000000000110101001110001; // input=2.552734375, output=-0.831575346677
			11'd654: out = 32'b10000000000000000110101010111000; // input=2.556640625, output=-0.833738574711
			11'd655: out = 32'b10000000000000000110101011111110; // input=2.560546875, output=-0.83588908092
			11'd656: out = 32'b10000000000000000110101101000100; // input=2.564453125, output=-0.83802683249
			11'd657: out = 32'b10000000000000000110101110001010; // input=2.568359375, output=-0.840151796802
			11'd658: out = 32'b10000000000000000110101111001111; // input=2.572265625, output=-0.842263941431
			11'd659: out = 32'b10000000000000000110110000010100; // input=2.576171875, output=-0.844363234149
			11'd660: out = 32'b10000000000000000110110001011000; // input=2.580078125, output=-0.846449642922
			11'd661: out = 32'b10000000000000000110110010011100; // input=2.583984375, output=-0.848523135916
			11'd662: out = 32'b10000000000000000110110011100000; // input=2.587890625, output=-0.85058368149
			11'd663: out = 32'b10000000000000000110110100100011; // input=2.591796875, output=-0.852631248204
			11'd664: out = 32'b10000000000000000110110101100110; // input=2.595703125, output=-0.854665804814
			11'd665: out = 32'b10000000000000000110110110101000; // input=2.599609375, output=-0.856687320275
			11'd666: out = 32'b10000000000000000110110111101010; // input=2.603515625, output=-0.858695763742
			11'd667: out = 32'b10000000000000000110111000101011; // input=2.607421875, output=-0.860691104568
			11'd668: out = 32'b10000000000000000110111001101100; // input=2.611328125, output=-0.862673312307
			11'd669: out = 32'b10000000000000000110111010101101; // input=2.615234375, output=-0.864642356712
			11'd670: out = 32'b10000000000000000110111011101101; // input=2.619140625, output=-0.866598207739
			11'd671: out = 32'b10000000000000000110111100101100; // input=2.623046875, output=-0.868540835543
			11'd672: out = 32'b10000000000000000110111101101100; // input=2.626953125, output=-0.870470210483
			11'd673: out = 32'b10000000000000000110111110101010; // input=2.630859375, output=-0.872386303118
			11'd674: out = 32'b10000000000000000110111111101001; // input=2.634765625, output=-0.874289084212
			11'd675: out = 32'b10000000000000000111000000100111; // input=2.638671875, output=-0.87617852473
			11'd676: out = 32'b10000000000000000111000001100100; // input=2.642578125, output=-0.878054595842
			11'd677: out = 32'b10000000000000000111000010100001; // input=2.646484375, output=-0.879917268921
			11'd678: out = 32'b10000000000000000111000011011110; // input=2.650390625, output=-0.881766515544
			11'd679: out = 32'b10000000000000000111000100011010; // input=2.654296875, output=-0.883602307496
			11'd680: out = 32'b10000000000000000111000101010110; // input=2.658203125, output=-0.885424616764
			11'd681: out = 32'b10000000000000000111000110010001; // input=2.662109375, output=-0.887233415541
			11'd682: out = 32'b10000000000000000111000111001100; // input=2.666015625, output=-0.889028676228
			11'd683: out = 32'b10000000000000000111001000000110; // input=2.669921875, output=-0.890810371432
			11'd684: out = 32'b10000000000000000111001001000000; // input=2.673828125, output=-0.892578473965
			11'd685: out = 32'b10000000000000000111001001111010; // input=2.677734375, output=-0.894332956848
			11'd686: out = 32'b10000000000000000111001010110011; // input=2.681640625, output=-0.896073793311
			11'd687: out = 32'b10000000000000000111001011101011; // input=2.685546875, output=-0.897800956791
			11'd688: out = 32'b10000000000000000111001100100011; // input=2.689453125, output=-0.899514420932
			11'd689: out = 32'b10000000000000000111001101011011; // input=2.693359375, output=-0.90121415959
			11'd690: out = 32'b10000000000000000111001110010010; // input=2.697265625, output=-0.902900146829
			11'd691: out = 32'b10000000000000000111001111001001; // input=2.701171875, output=-0.904572356923
			11'd692: out = 32'b10000000000000000111001111111111; // input=2.705078125, output=-0.906230764355
			11'd693: out = 32'b10000000000000000111010000110101; // input=2.708984375, output=-0.907875343821
			11'd694: out = 32'b10000000000000000111010001101011; // input=2.712890625, output=-0.909506070226
			11'd695: out = 32'b10000000000000000111010010100000; // input=2.716796875, output=-0.911122918687
			11'd696: out = 32'b10000000000000000111010011010100; // input=2.720703125, output=-0.912725864533
			11'd697: out = 32'b10000000000000000111010100001000; // input=2.724609375, output=-0.914314883306
			11'd698: out = 32'b10000000000000000111010100111100; // input=2.728515625, output=-0.915889950759
			11'd699: out = 32'b10000000000000000111010101101111; // input=2.732421875, output=-0.917451042858
			11'd700: out = 32'b10000000000000000111010110100010; // input=2.736328125, output=-0.918998135783
			11'd701: out = 32'b10000000000000000111010111010100; // input=2.740234375, output=-0.920531205927
			11'd702: out = 32'b10000000000000000111011000000110; // input=2.744140625, output=-0.922050229897
			11'd703: out = 32'b10000000000000000111011000110111; // input=2.748046875, output=-0.923555184515
			11'd704: out = 32'b10000000000000000111011001101000; // input=2.751953125, output=-0.925046046817
			11'd705: out = 32'b10000000000000000111011010011000; // input=2.755859375, output=-0.926522794055
			11'd706: out = 32'b10000000000000000111011011001000; // input=2.759765625, output=-0.927985403695
			11'd707: out = 32'b10000000000000000111011011111000; // input=2.763671875, output=-0.929433853419
			11'd708: out = 32'b10000000000000000111011100100111; // input=2.767578125, output=-0.930868121127
			11'd709: out = 32'b10000000000000000111011101010101; // input=2.771484375, output=-0.932288184932
			11'd710: out = 32'b10000000000000000111011110000011; // input=2.775390625, output=-0.933694023166
			11'd711: out = 32'b10000000000000000111011110110001; // input=2.779296875, output=-0.935085614378
			11'd712: out = 32'b10000000000000000111011111011110; // input=2.783203125, output=-0.936462937335
			11'd713: out = 32'b10000000000000000111100000001011; // input=2.787109375, output=-0.937825971019
			11'd714: out = 32'b10000000000000000111100000110111; // input=2.791015625, output=-0.939174694632
			11'd715: out = 32'b10000000000000000111100001100011; // input=2.794921875, output=-0.940509087596
			11'd716: out = 32'b10000000000000000111100010001110; // input=2.798828125, output=-0.941829129547
			11'd717: out = 32'b10000000000000000111100010111001; // input=2.802734375, output=-0.943134800345
			11'd718: out = 32'b10000000000000000111100011100011; // input=2.806640625, output=-0.944426080067
			11'd719: out = 32'b10000000000000000111100100001101; // input=2.810546875, output=-0.945702949008
			11'd720: out = 32'b10000000000000000111100100110110; // input=2.814453125, output=-0.946965387686
			11'd721: out = 32'b10000000000000000111100101011111; // input=2.818359375, output=-0.948213376837
			11'd722: out = 32'b10000000000000000111100110000111; // input=2.822265625, output=-0.949446897419
			11'd723: out = 32'b10000000000000000111100110101111; // input=2.826171875, output=-0.950665930609
			11'd724: out = 32'b10000000000000000111100111010111; // input=2.830078125, output=-0.951870457806
			11'd725: out = 32'b10000000000000000111100111111110; // input=2.833984375, output=-0.953060460632
			11'd726: out = 32'b10000000000000000111101000100100; // input=2.837890625, output=-0.954235920927
			11'd727: out = 32'b10000000000000000111101001001010; // input=2.841796875, output=-0.955396820757
			11'd728: out = 32'b10000000000000000111101001110000; // input=2.845703125, output=-0.956543142406
			11'd729: out = 32'b10000000000000000111101010010101; // input=2.849609375, output=-0.957674868384
			11'd730: out = 32'b10000000000000000111101010111010; // input=2.853515625, output=-0.958791981422
			11'd731: out = 32'b10000000000000000111101011011110; // input=2.857421875, output=-0.959894464473
			11'd732: out = 32'b10000000000000000111101100000001; // input=2.861328125, output=-0.960982300717
			11'd733: out = 32'b10000000000000000111101100100101; // input=2.865234375, output=-0.962055473552
			11'd734: out = 32'b10000000000000000111101101000111; // input=2.869140625, output=-0.963113966605
			11'd735: out = 32'b10000000000000000111101101101010; // input=2.873046875, output=-0.964157763723
			11'd736: out = 32'b10000000000000000111101110001011; // input=2.876953125, output=-0.965186848981
			11'd737: out = 32'b10000000000000000111101110101100; // input=2.880859375, output=-0.966201206674
			11'd738: out = 32'b10000000000000000111101111001101; // input=2.884765625, output=-0.967200821326
			11'd739: out = 32'b10000000000000000111101111101110; // input=2.888671875, output=-0.968185677683
			11'd740: out = 32'b10000000000000000111110000001101; // input=2.892578125, output=-0.969155760718
			11'd741: out = 32'b10000000000000000111110000101101; // input=2.896484375, output=-0.970111055629
			11'd742: out = 32'b10000000000000000111110001001011; // input=2.900390625, output=-0.971051547838
			11'd743: out = 32'b10000000000000000111110001101010; // input=2.904296875, output=-0.971977222996
			11'd744: out = 32'b10000000000000000111110010001000; // input=2.908203125, output=-0.972888066977
			11'd745: out = 32'b10000000000000000111110010100101; // input=2.912109375, output=-0.973784065883
			11'd746: out = 32'b10000000000000000111110011000010; // input=2.916015625, output=-0.974665206042
			11'd747: out = 32'b10000000000000000111110011011110; // input=2.919921875, output=-0.975531474009
			11'd748: out = 32'b10000000000000000111110011111010; // input=2.923828125, output=-0.976382856567
			11'd749: out = 32'b10000000000000000111110100010110; // input=2.927734375, output=-0.977219340723
			11'd750: out = 32'b10000000000000000111110100110000; // input=2.931640625, output=-0.978040913714
			11'd751: out = 32'b10000000000000000111110101001011; // input=2.935546875, output=-0.978847563005
			11'd752: out = 32'b10000000000000000111110101100101; // input=2.939453125, output=-0.979639276285
			11'd753: out = 32'b10000000000000000111110101111110; // input=2.943359375, output=-0.980416041476
			11'd754: out = 32'b10000000000000000111110110010111; // input=2.947265625, output=-0.981177846724
			11'd755: out = 32'b10000000000000000111110110110000; // input=2.951171875, output=-0.981924680406
			11'd756: out = 32'b10000000000000000111110111001000; // input=2.955078125, output=-0.982656531125
			11'd757: out = 32'b10000000000000000111110111011111; // input=2.958984375, output=-0.983373387714
			11'd758: out = 32'b10000000000000000111110111110110; // input=2.962890625, output=-0.984075239235
			11'd759: out = 32'b10000000000000000111111000001101; // input=2.966796875, output=-0.984762074979
			11'd760: out = 32'b10000000000000000111111000100011; // input=2.970703125, output=-0.985433884466
			11'd761: out = 32'b10000000000000000111111000111000; // input=2.974609375, output=-0.986090657443
			11'd762: out = 32'b10000000000000000111111001001101; // input=2.978515625, output=-0.986732383891
			11'd763: out = 32'b10000000000000000111111001100010; // input=2.982421875, output=-0.987359054016
			11'd764: out = 32'b10000000000000000111111001110110; // input=2.986328125, output=-0.987970658257
			11'd765: out = 32'b10000000000000000111111010001001; // input=2.990234375, output=-0.988567187281
			11'd766: out = 32'b10000000000000000111111010011100; // input=2.994140625, output=-0.989148631986
			11'd767: out = 32'b10000000000000000111111010101111; // input=2.998046875, output=-0.9897149835
			11'd768: out = 32'b10000000000000000111111011000001; // input=3.001953125, output=-0.990266233181
			11'd769: out = 32'b10000000000000000111111011010011; // input=3.005859375, output=-0.990802372617
			11'd770: out = 32'b10000000000000000111111011100100; // input=3.009765625, output=-0.991323393629
			11'd771: out = 32'b10000000000000000111111011110100; // input=3.013671875, output=-0.991829288265
			11'd772: out = 32'b10000000000000000111111100000100; // input=3.017578125, output=-0.992320048806
			11'd773: out = 32'b10000000000000000111111100010100; // input=3.021484375, output=-0.992795667765
			11'd774: out = 32'b10000000000000000111111100100011; // input=3.025390625, output=-0.993256137883
			11'd775: out = 32'b10000000000000000111111100110010; // input=3.029296875, output=-0.993701452134
			11'd776: out = 32'b10000000000000000111111101000000; // input=3.033203125, output=-0.994131603724
			11'd777: out = 32'b10000000000000000111111101001101; // input=3.037109375, output=-0.994546586089
			11'd778: out = 32'b10000000000000000111111101011010; // input=3.041015625, output=-0.994946392896
			11'd779: out = 32'b10000000000000000111111101100111; // input=3.044921875, output=-0.995331018046
			11'd780: out = 32'b10000000000000000111111101110011; // input=3.048828125, output=-0.995700455669
			11'd781: out = 32'b10000000000000000111111101111111; // input=3.052734375, output=-0.996054700128
			11'd782: out = 32'b10000000000000000111111110001010; // input=3.056640625, output=-0.996393746017
			11'd783: out = 32'b10000000000000000111111110010100; // input=3.060546875, output=-0.996717588164
			11'd784: out = 32'b10000000000000000111111110011111; // input=3.064453125, output=-0.997026221627
			11'd785: out = 32'b10000000000000000111111110101000; // input=3.068359375, output=-0.997319641697
			11'd786: out = 32'b10000000000000000111111110110001; // input=3.072265625, output=-0.997597843896
			11'd787: out = 32'b10000000000000000111111110111010; // input=3.076171875, output=-0.997860823979
			11'd788: out = 32'b10000000000000000111111111000010; // input=3.080078125, output=-0.998108577933
			11'd789: out = 32'b10000000000000000111111111001010; // input=3.083984375, output=-0.998341101979
			11'd790: out = 32'b10000000000000000111111111010001; // input=3.087890625, output=-0.998558392568
			11'd791: out = 32'b10000000000000000111111111010111; // input=3.091796875, output=-0.998760446384
			11'd792: out = 32'b10000000000000000111111111011110; // input=3.095703125, output=-0.998947260345
			11'd793: out = 32'b10000000000000000111111111100011; // input=3.099609375, output=-0.999118831599
			11'd794: out = 32'b10000000000000000111111111101000; // input=3.103515625, output=-0.99927515753
			11'd795: out = 32'b10000000000000000111111111101101; // input=3.107421875, output=-0.999416235751
			11'd796: out = 32'b10000000000000000111111111110001; // input=3.111328125, output=-0.99954206411
			11'd797: out = 32'b10000000000000000111111111110101; // input=3.115234375, output=-0.999652640687
			11'd798: out = 32'b10000000000000000111111111111000; // input=3.119140625, output=-0.999747963794
			11'd799: out = 32'b10000000000000000111111111111010; // input=3.123046875, output=-0.999828031977
			11'd800: out = 32'b10000000000000000111111111111100; // input=3.126953125, output=-0.999892844015
			11'd801: out = 32'b10000000000000000111111111111110; // input=3.130859375, output=-0.999942398918
			11'd802: out = 32'b10000000000000000111111111111111; // input=3.134765625, output=-0.999976695931
			11'd803: out = 32'b10000000000000000111111111111111; // input=3.138671875, output=-0.999995734529
			11'd804: out = 32'b10000000000000000111111111111111; // input=3.142578125, output=-0.999999514423
			11'd805: out = 32'b10000000000000000111111111111111; // input=3.146484375, output=-0.999988035555
			11'd806: out = 32'b10000000000000000111111111111111; // input=3.150390625, output=-0.999961298099
			11'd807: out = 32'b10000000000000000111111111111101; // input=3.154296875, output=-0.999919302465
			11'd808: out = 32'b10000000000000000111111111111011; // input=3.158203125, output=-0.999862049292
			11'd809: out = 32'b10000000000000000111111111111001; // input=3.162109375, output=-0.999789539454
			11'd810: out = 32'b10000000000000000111111111110110; // input=3.166015625, output=-0.999701774058
			11'd811: out = 32'b10000000000000000111111111110011; // input=3.169921875, output=-0.999598754443
			11'd812: out = 32'b10000000000000000111111111101111; // input=3.173828125, output=-0.999480482181
			11'd813: out = 32'b10000000000000000111111111101011; // input=3.177734375, output=-0.999346959076
			11'd814: out = 32'b10000000000000000111111111100110; // input=3.181640625, output=-0.999198187167
			11'd815: out = 32'b10000000000000000111111111100000; // input=3.185546875, output=-0.999034168722
			11'd816: out = 32'b10000000000000000111111111011010; // input=3.189453125, output=-0.998854906245
			11'd817: out = 32'b10000000000000000111111111010100; // input=3.193359375, output=-0.998660402471
			11'd818: out = 32'b10000000000000000111111111001101; // input=3.197265625, output=-0.998450660368
			11'd819: out = 32'b10000000000000000111111111000110; // input=3.201171875, output=-0.998225683137
			11'd820: out = 32'b10000000000000000111111110111110; // input=3.205078125, output=-0.997985474209
			11'd821: out = 32'b10000000000000000111111110110110; // input=3.208984375, output=-0.997730037251
			11'd822: out = 32'b10000000000000000111111110101101; // input=3.212890625, output=-0.997459376161
			11'd823: out = 32'b10000000000000000111111110100011; // input=3.216796875, output=-0.997173495067
			11'd824: out = 32'b10000000000000000111111110011010; // input=3.220703125, output=-0.996872398333
			11'd825: out = 32'b10000000000000000111111110001111; // input=3.224609375, output=-0.996556090553
			11'd826: out = 32'b10000000000000000111111110000100; // input=3.228515625, output=-0.996224576552
			11'd827: out = 32'b10000000000000000111111101111001; // input=3.232421875, output=-0.995877861391
			11'd828: out = 32'b10000000000000000111111101101101; // input=3.236328125, output=-0.995515950358
			11'd829: out = 32'b10000000000000000111111101100001; // input=3.240234375, output=-0.995138848977
			11'd830: out = 32'b10000000000000000111111101010100; // input=3.244140625, output=-0.994746563001
			11'd831: out = 32'b10000000000000000111111101000111; // input=3.248046875, output=-0.994339098417
			11'd832: out = 32'b10000000000000000111111100111001; // input=3.251953125, output=-0.993916461441
			11'd833: out = 32'b10000000000000000111111100101010; // input=3.255859375, output=-0.993478658524
			11'd834: out = 32'b10000000000000000111111100011011; // input=3.259765625, output=-0.993025696344
			11'd835: out = 32'b10000000000000000111111100001100; // input=3.263671875, output=-0.992557581813
			11'd836: out = 32'b10000000000000000111111011111100; // input=3.267578125, output=-0.992074322076
			11'd837: out = 32'b10000000000000000111111011101100; // input=3.271484375, output=-0.991575924504
			11'd838: out = 32'b10000000000000000111111011011011; // input=3.275390625, output=-0.991062396704
			11'd839: out = 32'b10000000000000000111111011001010; // input=3.279296875, output=-0.990533746511
			11'd840: out = 32'b10000000000000000111111010111000; // input=3.283203125, output=-0.989989981992
			11'd841: out = 32'b10000000000000000111111010100110; // input=3.287109375, output=-0.989431111444
			11'd842: out = 32'b10000000000000000111111010010011; // input=3.291015625, output=-0.988857143395
			11'd843: out = 32'b10000000000000000111111010000000; // input=3.294921875, output=-0.988268086602
			11'd844: out = 32'b10000000000000000111111001101100; // input=3.298828125, output=-0.987663950053
			11'd845: out = 32'b10000000000000000111111001010111; // input=3.302734375, output=-0.987044742969
			11'd846: out = 32'b10000000000000000111111001000011; // input=3.306640625, output=-0.986410474795
			11'd847: out = 32'b10000000000000000111111000101101; // input=3.310546875, output=-0.985761155212
			11'd848: out = 32'b10000000000000000111111000011000; // input=3.314453125, output=-0.985096794126
			11'd849: out = 32'b10000000000000000111111000000001; // input=3.318359375, output=-0.984417401675
			11'd850: out = 32'b10000000000000000111110111101011; // input=3.322265625, output=-0.983722988226
			11'd851: out = 32'b10000000000000000111110111010011; // input=3.326171875, output=-0.983013564374
			11'd852: out = 32'b10000000000000000111110110111100; // input=3.330078125, output=-0.982289140945
			11'd853: out = 32'b10000000000000000111110110100011; // input=3.333984375, output=-0.981549728992
			11'd854: out = 32'b10000000000000000111110110001011; // input=3.337890625, output=-0.980795339798
			11'd855: out = 32'b10000000000000000111110101110001; // input=3.341796875, output=-0.980025984873
			11'd856: out = 32'b10000000000000000111110101011000; // input=3.345703125, output=-0.979241675958
			11'd857: out = 32'b10000000000000000111110100111110; // input=3.349609375, output=-0.978442425019
			11'd858: out = 32'b10000000000000000111110100100011; // input=3.353515625, output=-0.977628244254
			11'd859: out = 32'b10000000000000000111110100001000; // input=3.357421875, output=-0.976799146083
			11'd860: out = 32'b10000000000000000111110011101100; // input=3.361328125, output=-0.97595514316
			11'd861: out = 32'b10000000000000000111110011010000; // input=3.365234375, output=-0.975096248362
			11'd862: out = 32'b10000000000000000111110010110011; // input=3.369140625, output=-0.974222474795
			11'd863: out = 32'b10000000000000000111110010010110; // input=3.373046875, output=-0.973333835791
			11'd864: out = 32'b10000000000000000111110001111001; // input=3.376953125, output=-0.972430344911
			11'd865: out = 32'b10000000000000000111110001011011; // input=3.380859375, output=-0.97151201594
			11'd866: out = 32'b10000000000000000111110000111100; // input=3.384765625, output=-0.970578862891
			11'd867: out = 32'b10000000000000000111110000011101; // input=3.388671875, output=-0.969630900003
			11'd868: out = 32'b10000000000000000111101111111101; // input=3.392578125, output=-0.96866814174
			11'd869: out = 32'b10000000000000000111101111011101; // input=3.396484375, output=-0.967690602793
			11'd870: out = 32'b10000000000000000111101110111101; // input=3.400390625, output=-0.966698298078
			11'd871: out = 32'b10000000000000000111101110011100; // input=3.404296875, output=-0.965691242737
			11'd872: out = 32'b10000000000000000111101101111010; // input=3.408203125, output=-0.964669452135
			11'd873: out = 32'b10000000000000000111101101011000; // input=3.412109375, output=-0.963632941864
			11'd874: out = 32'b10000000000000000111101100110110; // input=3.416015625, output=-0.96258172774
			11'd875: out = 32'b10000000000000000111101100010011; // input=3.419921875, output=-0.961515825803
			11'd876: out = 32'b10000000000000000111101011110000; // input=3.423828125, output=-0.960435252318
			11'd877: out = 32'b10000000000000000111101011001100; // input=3.427734375, output=-0.959340023773
			11'd878: out = 32'b10000000000000000111101010100111; // input=3.431640625, output=-0.958230156879
			11'd879: out = 32'b10000000000000000111101010000010; // input=3.435546875, output=-0.957105668571
			11'd880: out = 32'b10000000000000000111101001011101; // input=3.439453125, output=-0.955966576009
			11'd881: out = 32'b10000000000000000111101000110111; // input=3.443359375, output=-0.954812896573
			11'd882: out = 32'b10000000000000000111101000010001; // input=3.447265625, output=-0.953644647867
			11'd883: out = 32'b10000000000000000111100111101010; // input=3.451171875, output=-0.952461847717
			11'd884: out = 32'b10000000000000000111100111000011; // input=3.455078125, output=-0.951264514171
			11'd885: out = 32'b10000000000000000111100110011011; // input=3.458984375, output=-0.950052665499
			11'd886: out = 32'b10000000000000000111100101110011; // input=3.462890625, output=-0.948826320192
			11'd887: out = 32'b10000000000000000111100101001010; // input=3.466796875, output=-0.947585496963
			11'd888: out = 32'b10000000000000000111100100100001; // input=3.470703125, output=-0.946330214745
			11'd889: out = 32'b10000000000000000111100011111000; // input=3.474609375, output=-0.945060492692
			11'd890: out = 32'b10000000000000000111100011001110; // input=3.478515625, output=-0.943776350179
			11'd891: out = 32'b10000000000000000111100010100011; // input=3.482421875, output=-0.9424778068
			11'd892: out = 32'b10000000000000000111100001111000; // input=3.486328125, output=-0.94116488237
			11'd893: out = 32'b10000000000000000111100001001101; // input=3.490234375, output=-0.939837596921
			11'd894: out = 32'b10000000000000000111100000100001; // input=3.494140625, output=-0.938495970706
			11'd895: out = 32'b10000000000000000111011111110100; // input=3.498046875, output=-0.937140024198
			11'd896: out = 32'b10000000000000000111011111000111; // input=3.501953125, output=-0.935769778086
			11'd897: out = 32'b10000000000000000111011110011010; // input=3.505859375, output=-0.934385253279
			11'd898: out = 32'b10000000000000000111011101101100; // input=3.509765625, output=-0.932986470902
			11'd899: out = 32'b10000000000000000111011100111110; // input=3.513671875, output=-0.931573452299
			11'd900: out = 32'b10000000000000000111011100001111; // input=3.517578125, output=-0.930146219032
			11'd901: out = 32'b10000000000000000111011011100000; // input=3.521484375, output=-0.928704792878
			11'd902: out = 32'b10000000000000000111011010110000; // input=3.525390625, output=-0.927249195831
			11'd903: out = 32'b10000000000000000111011010000000; // input=3.529296875, output=-0.925779450103
			11'd904: out = 32'b10000000000000000111011001001111; // input=3.533203125, output=-0.924295578119
			11'd905: out = 32'b10000000000000000111011000011110; // input=3.537109375, output=-0.922797602521
			11'd906: out = 32'b10000000000000000111010111101101; // input=3.541015625, output=-0.921285546168
			11'd907: out = 32'b10000000000000000111010110111011; // input=3.544921875, output=-0.919759432131
			11'd908: out = 32'b10000000000000000111010110001000; // input=3.548828125, output=-0.918219283696
			11'd909: out = 32'b10000000000000000111010101010101; // input=3.552734375, output=-0.916665124365
			11'd910: out = 32'b10000000000000000111010100100010; // input=3.556640625, output=-0.915096977852
			11'd911: out = 32'b10000000000000000111010011101110; // input=3.560546875, output=-0.913514868085
			11'd912: out = 32'b10000000000000000111010010111010; // input=3.564453125, output=-0.911918819205
			11'd913: out = 32'b10000000000000000111010010000101; // input=3.568359375, output=-0.910308855566
			11'd914: out = 32'b10000000000000000111010001010000; // input=3.572265625, output=-0.908685001733
			11'd915: out = 32'b10000000000000000111010000011010; // input=3.576171875, output=-0.907047282486
			11'd916: out = 32'b10000000000000000111001111100100; // input=3.580078125, output=-0.905395722813
			11'd917: out = 32'b10000000000000000111001110101101; // input=3.583984375, output=-0.903730347915
			11'd918: out = 32'b10000000000000000111001101110110; // input=3.587890625, output=-0.902051183204
			11'd919: out = 32'b10000000000000000111001100111111; // input=3.591796875, output=-0.900358254301
			11'd920: out = 32'b10000000000000000111001100000111; // input=3.595703125, output=-0.89865158704
			11'd921: out = 32'b10000000000000000111001011001111; // input=3.599609375, output=-0.896931207461
			11'd922: out = 32'b10000000000000000111001010010110; // input=3.603515625, output=-0.895197141815
			11'd923: out = 32'b10000000000000000111001001011101; // input=3.607421875, output=-0.893449416562
			11'd924: out = 32'b10000000000000000111001000100011; // input=3.611328125, output=-0.89168805837
			11'd925: out = 32'b10000000000000000111000111101001; // input=3.615234375, output=-0.889913094116
			11'd926: out = 32'b10000000000000000111000110101110; // input=3.619140625, output=-0.888124550883
			11'd927: out = 32'b10000000000000000111000101110011; // input=3.623046875, output=-0.886322455962
			11'd928: out = 32'b10000000000000000111000100111000; // input=3.626953125, output=-0.88450683685
			11'd929: out = 32'b10000000000000000111000011111100; // input=3.630859375, output=-0.882677721253
			11'd930: out = 32'b10000000000000000111000010111111; // input=3.634765625, output=-0.880835137079
			11'd931: out = 32'b10000000000000000111000010000010; // input=3.638671875, output=-0.878979112445
			11'd932: out = 32'b10000000000000000111000001000101; // input=3.642578125, output=-0.877109675671
			11'd933: out = 32'b10000000000000000111000000000111; // input=3.646484375, output=-0.875226855283
			11'd934: out = 32'b10000000000000000110111111001001; // input=3.650390625, output=-0.87333068001
			11'd935: out = 32'b10000000000000000110111110001011; // input=3.654296875, output=-0.871421178785
			11'd936: out = 32'b10000000000000000110111101001100; // input=3.658203125, output=-0.869498380745
			11'd937: out = 32'b10000000000000000110111100001100; // input=3.662109375, output=-0.867562315229
			11'd938: out = 32'b10000000000000000110111011001100; // input=3.666015625, output=-0.86561301178
			11'd939: out = 32'b10000000000000000110111010001100; // input=3.669921875, output=-0.863650500142
			11'd940: out = 32'b10000000000000000110111001001011; // input=3.673828125, output=-0.861674810259
			11'd941: out = 32'b10000000000000000110111000001010; // input=3.677734375, output=-0.859685972279
			11'd942: out = 32'b10000000000000000110110111001001; // input=3.681640625, output=-0.857684016548
			11'd943: out = 32'b10000000000000000110110110000111; // input=3.685546875, output=-0.855668973615
			11'd944: out = 32'b10000000000000000110110101000100; // input=3.689453125, output=-0.853640874226
			11'd945: out = 32'b10000000000000000110110100000001; // input=3.693359375, output=-0.851599749328
			11'd946: out = 32'b10000000000000000110110010111110; // input=3.697265625, output=-0.849545630065
			11'd947: out = 32'b10000000000000000110110001111010; // input=3.701171875, output=-0.847478547781
			11'd948: out = 32'b10000000000000000110110000110110; // input=3.705078125, output=-0.845398534017
			11'd949: out = 32'b10000000000000000110101111110001; // input=3.708984375, output=-0.843305620512
			11'd950: out = 32'b10000000000000000110101110101100; // input=3.712890625, output=-0.8411998392
			11'd951: out = 32'b10000000000000000110101101100111; // input=3.716796875, output=-0.839081222214
			11'd952: out = 32'b10000000000000000110101100100001; // input=3.720703125, output=-0.83694980188
			11'd953: out = 32'b10000000000000000110101011011011; // input=3.724609375, output=-0.834805610723
			11'd954: out = 32'b10000000000000000110101010010100; // input=3.728515625, output=-0.832648681459
			11'd955: out = 32'b10000000000000000110101001001101; // input=3.732421875, output=-0.830479047
			11'd956: out = 32'b10000000000000000110101000000110; // input=3.736328125, output=-0.828296740453
			11'd957: out = 32'b10000000000000000110100110111110; // input=3.740234375, output=-0.826101795117
			11'd958: out = 32'b10000000000000000110100101110101; // input=3.744140625, output=-0.823894244484
			11'd959: out = 32'b10000000000000000110100100101101; // input=3.748046875, output=-0.821674122238
			11'd960: out = 32'b10000000000000000110100011100011; // input=3.751953125, output=-0.819441462256
			11'd961: out = 32'b10000000000000000110100010011010; // input=3.755859375, output=-0.817196298606
			11'd962: out = 32'b10000000000000000110100001010000; // input=3.759765625, output=-0.814938665546
			11'd963: out = 32'b10000000000000000110100000000110; // input=3.763671875, output=-0.812668597524
			11'd964: out = 32'b10000000000000000110011110111011; // input=3.767578125, output=-0.810386129179
			11'd965: out = 32'b10000000000000000110011101110000; // input=3.771484375, output=-0.808091295339
			11'd966: out = 32'b10000000000000000110011100100100; // input=3.775390625, output=-0.80578413102
			11'd967: out = 32'b10000000000000000110011011011000; // input=3.779296875, output=-0.803464671426
			11'd968: out = 32'b10000000000000000110011010001100; // input=3.783203125, output=-0.801132951951
			11'd969: out = 32'b10000000000000000110011000111111; // input=3.787109375, output=-0.798789008172
			11'd970: out = 32'b10000000000000000110010111110010; // input=3.791015625, output=-0.796432875855
			11'd971: out = 32'b10000000000000000110010110100100; // input=3.794921875, output=-0.794064590953
			11'd972: out = 32'b10000000000000000110010101010110; // input=3.798828125, output=-0.791684189602
			11'd973: out = 32'b10000000000000000110010100001000; // input=3.802734375, output=-0.789291708124
			11'd974: out = 32'b10000000000000000110010010111001; // input=3.806640625, output=-0.786887183026
			11'd975: out = 32'b10000000000000000110010001101010; // input=3.810546875, output=-0.784470650998
			11'd976: out = 32'b10000000000000000110010000011010; // input=3.814453125, output=-0.782042148913
			11'd977: out = 32'b10000000000000000110001111001010; // input=3.818359375, output=-0.779601713826
			11'd978: out = 32'b10000000000000000110001101111010; // input=3.822265625, output=-0.777149382977
			11'd979: out = 32'b10000000000000000110001100101001; // input=3.826171875, output=-0.774685193784
			11'd980: out = 32'b10000000000000000110001011011000; // input=3.830078125, output=-0.772209183849
			11'd981: out = 32'b10000000000000000110001010000110; // input=3.833984375, output=-0.769721390951
			11'd982: out = 32'b10000000000000000110001000110100; // input=3.837890625, output=-0.767221853052
			11'd983: out = 32'b10000000000000000110000111100010; // input=3.841796875, output=-0.764710608291
			11'd984: out = 32'b10000000000000000110000110001111; // input=3.845703125, output=-0.762187694988
			11'd985: out = 32'b10000000000000000110000100111100; // input=3.849609375, output=-0.759653151638
			11'd986: out = 32'b10000000000000000110000011101001; // input=3.853515625, output=-0.757107016915
			11'd987: out = 32'b10000000000000000110000010010101; // input=3.857421875, output=-0.754549329671
			11'd988: out = 32'b10000000000000000110000001000001; // input=3.861328125, output=-0.751980128932
			11'd989: out = 32'b10000000000000000101111111101100; // input=3.865234375, output=-0.749399453902
			11'd990: out = 32'b10000000000000000101111110010111; // input=3.869140625, output=-0.746807343958
			11'd991: out = 32'b10000000000000000101111101000010; // input=3.873046875, output=-0.744203838653
			11'd992: out = 32'b10000000000000000101111011101100; // input=3.876953125, output=-0.741588977713
			11'd993: out = 32'b10000000000000000101111010010110; // input=3.880859375, output=-0.738962801038
			11'd994: out = 32'b10000000000000000101111001000000; // input=3.884765625, output=-0.736325348699
			11'd995: out = 32'b10000000000000000101110111101001; // input=3.888671875, output=-0.733676660942
			11'd996: out = 32'b10000000000000000101110110010010; // input=3.892578125, output=-0.731016778181
			11'd997: out = 32'b10000000000000000101110100111010; // input=3.896484375, output=-0.728345741004
			11'd998: out = 32'b10000000000000000101110011100011; // input=3.900390625, output=-0.725663590167
			11'd999: out = 32'b10000000000000000101110010001010; // input=3.904296875, output=-0.722970366596
			11'd1000: out = 32'b10000000000000000101110000110010; // input=3.908203125, output=-0.720266111387
			11'd1001: out = 32'b10000000000000000101101111011001; // input=3.912109375, output=-0.717550865803
			11'd1002: out = 32'b10000000000000000101101101111111; // input=3.916015625, output=-0.714824671276
			11'd1003: out = 32'b10000000000000000101101100100110; // input=3.919921875, output=-0.712087569404
			11'd1004: out = 32'b10000000000000000101101011001100; // input=3.923828125, output=-0.709339601952
			11'd1005: out = 32'b10000000000000000101101001110001; // input=3.927734375, output=-0.70658081085
			11'd1006: out = 32'b10000000000000000101101000010110; // input=3.931640625, output=-0.703811238194
			11'd1007: out = 32'b10000000000000000101100110111011; // input=3.935546875, output=-0.701030926245
			11'd1008: out = 32'b10000000000000000101100101100000; // input=3.939453125, output=-0.698239917426
			11'd1009: out = 32'b10000000000000000101100100000100; // input=3.943359375, output=-0.695438254325
			11'd1010: out = 32'b10000000000000000101100010101000; // input=3.947265625, output=-0.692625979692
			11'd1011: out = 32'b10000000000000000101100001001011; // input=3.951171875, output=-0.689803136439
			11'd1012: out = 32'b10000000000000000101011111101111; // input=3.955078125, output=-0.686969767639
			11'd1013: out = 32'b10000000000000000101011110010001; // input=3.958984375, output=-0.684125916525
			11'd1014: out = 32'b10000000000000000101011100110100; // input=3.962890625, output=-0.681271626491
			11'd1015: out = 32'b10000000000000000101011011010110; // input=3.966796875, output=-0.678406941091
			11'd1016: out = 32'b10000000000000000101011001111000; // input=3.970703125, output=-0.675531904035
			11'd1017: out = 32'b10000000000000000101011000011001; // input=3.974609375, output=-0.672646559194
			11'd1018: out = 32'b10000000000000000101010110111010; // input=3.978515625, output=-0.669750950593
			11'd1019: out = 32'b10000000000000000101010101011011; // input=3.982421875, output=-0.666845122418
			11'd1020: out = 32'b10000000000000000101010011111100; // input=3.986328125, output=-0.663929119006
			11'd1021: out = 32'b10000000000000000101010010011100; // input=3.990234375, output=-0.661002984852
			11'd1022: out = 32'b10000000000000000101010000111100; // input=3.994140625, output=-0.658066764607
			11'd1023: out = 32'b10000000000000000101001111011011; // input=3.998046875, output=-0.655120503072
			11'd1024: out = 32'b00000000000000000111111111111111; // input=-0.001953125, output=0.999998092652
			11'd1025: out = 32'b00000000000000000111111111111111; // input=-0.005859375, output=0.999982833911
			11'd1026: out = 32'b00000000000000000111111111111110; // input=-0.009765625, output=0.999952316663
			11'd1027: out = 32'b00000000000000000111111111111101; // input=-0.013671875, output=0.999906541373
			11'd1028: out = 32'b00000000000000000111111111111011; // input=-0.017578125, output=0.999845508739
			11'd1029: out = 32'b00000000000000000111111111111000; // input=-0.021484375, output=0.999769219693
			11'd1030: out = 32'b00000000000000000111111111110101; // input=-0.025390625, output=0.999677675398
			11'd1031: out = 32'b00000000000000000111111111110010; // input=-0.029296875, output=0.999570877252
			11'd1032: out = 32'b00000000000000000111111111101110; // input=-0.033203125, output=0.999448826885
			11'd1033: out = 32'b00000000000000000111111111101001; // input=-0.037109375, output=0.999311526157
			11'd1034: out = 32'b00000000000000000111111111100100; // input=-0.041015625, output=0.999158977166
			11'd1035: out = 32'b00000000000000000111111111011111; // input=-0.044921875, output=0.998991182238
			11'd1036: out = 32'b00000000000000000111111111011001; // input=-0.048828125, output=0.998808143933
			11'd1037: out = 32'b00000000000000000111111111010010; // input=-0.052734375, output=0.998609865045
			11'd1038: out = 32'b00000000000000000111111111001011; // input=-0.056640625, output=0.998396348599
			11'd1039: out = 32'b00000000000000000111111111000100; // input=-0.060546875, output=0.998167597854
			11'd1040: out = 32'b00000000000000000111111110111100; // input=-0.064453125, output=0.997923616299
			11'd1041: out = 32'b00000000000000000111111110110011; // input=-0.068359375, output=0.997664407657
			11'd1042: out = 32'b00000000000000000111111110101010; // input=-0.072265625, output=0.997389975884
			11'd1043: out = 32'b00000000000000000111111110100001; // input=-0.076171875, output=0.997100325166
			11'd1044: out = 32'b00000000000000000111111110010111; // input=-0.080078125, output=0.996795459925
			11'd1045: out = 32'b00000000000000000111111110001101; // input=-0.083984375, output=0.996475384812
			11'd1046: out = 32'b00000000000000000111111110000010; // input=-0.087890625, output=0.99614010471
			11'd1047: out = 32'b00000000000000000111111101110110; // input=-0.091796875, output=0.995789624735
			11'd1048: out = 32'b00000000000000000111111101101010; // input=-0.095703125, output=0.995423950236
			11'd1049: out = 32'b00000000000000000111111101011110; // input=-0.099609375, output=0.995043086793
			11'd1050: out = 32'b00000000000000000111111101010001; // input=-0.103515625, output=0.994647040216
			11'd1051: out = 32'b00000000000000000111111101000011; // input=-0.107421875, output=0.994235816549
			11'd1052: out = 32'b00000000000000000111111100110101; // input=-0.111328125, output=0.993809422066
			11'd1053: out = 32'b00000000000000000111111100100111; // input=-0.115234375, output=0.993367863275
			11'd1054: out = 32'b00000000000000000111111100011000; // input=-0.119140625, output=0.992911146912
			11'd1055: out = 32'b00000000000000000111111100001000; // input=-0.123046875, output=0.992439279947
			11'd1056: out = 32'b00000000000000000111111011111000; // input=-0.126953125, output=0.991952269579
			11'd1057: out = 32'b00000000000000000111111011101000; // input=-0.130859375, output=0.99145012324
			11'd1058: out = 32'b00000000000000000111111011010111; // input=-0.134765625, output=0.990932848592
			11'd1059: out = 32'b00000000000000000111111011000101; // input=-0.138671875, output=0.990400453528
			11'd1060: out = 32'b00000000000000000111111010110100; // input=-0.142578125, output=0.989852946172
			11'd1061: out = 32'b00000000000000000111111010100001; // input=-0.146484375, output=0.989290334878
			11'd1062: out = 32'b00000000000000000111111010001110; // input=-0.150390625, output=0.98871262823
			11'd1063: out = 32'b00000000000000000111111001111011; // input=-0.154296875, output=0.988119835044
			11'd1064: out = 32'b00000000000000000111111001100111; // input=-0.158203125, output=0.987511964365
			11'd1065: out = 32'b00000000000000000111111001010010; // input=-0.162109375, output=0.986889025468
			11'd1066: out = 32'b00000000000000000111111000111101; // input=-0.166015625, output=0.986251027859
			11'd1067: out = 32'b00000000000000000111111000101000; // input=-0.169921875, output=0.985597981273
			11'd1068: out = 32'b00000000000000000111111000010010; // input=-0.173828125, output=0.984929895674
			11'd1069: out = 32'b00000000000000000111110111111100; // input=-0.177734375, output=0.984246781257
			11'd1070: out = 32'b00000000000000000111110111100101; // input=-0.181640625, output=0.983548648445
			11'd1071: out = 32'b00000000000000000111110111001110; // input=-0.185546875, output=0.98283550789
			11'd1072: out = 32'b00000000000000000111110110110110; // input=-0.189453125, output=0.982107370475
			11'd1073: out = 32'b00000000000000000111110110011101; // input=-0.193359375, output=0.98136424731
			11'd1074: out = 32'b00000000000000000111110110000101; // input=-0.197265625, output=0.980606149734
			11'd1075: out = 32'b00000000000000000111110101101011; // input=-0.201171875, output=0.979833089314
			11'd1076: out = 32'b00000000000000000111110101010001; // input=-0.205078125, output=0.979045077847
			11'd1077: out = 32'b00000000000000000111110100110111; // input=-0.208984375, output=0.978242127357
			11'd1078: out = 32'b00000000000000000111110100011100; // input=-0.212890625, output=0.977424250095
			11'd1079: out = 32'b00000000000000000111110100000001; // input=-0.216796875, output=0.976591458542
			11'd1080: out = 32'b00000000000000000111110011100101; // input=-0.220703125, output=0.975743765405
			11'd1081: out = 32'b00000000000000000111110011001001; // input=-0.224609375, output=0.974881183619
			11'd1082: out = 32'b00000000000000000111110010101100; // input=-0.228515625, output=0.974003726345
			11'd1083: out = 32'b00000000000000000111110010001111; // input=-0.232421875, output=0.973111406972
			11'd1084: out = 32'b00000000000000000111110001110001; // input=-0.236328125, output=0.972204239117
			11'd1085: out = 32'b00000000000000000111110001010011; // input=-0.240234375, output=0.971282236621
			11'd1086: out = 32'b00000000000000000111110000110100; // input=-0.244140625, output=0.970345413553
			11'd1087: out = 32'b00000000000000000111110000010101; // input=-0.248046875, output=0.969393784208
			11'd1088: out = 32'b00000000000000000111101111110101; // input=-0.251953125, output=0.968427363107
			11'd1089: out = 32'b00000000000000000111101111010101; // input=-0.255859375, output=0.967446164995
			11'd1090: out = 32'b00000000000000000111101110110101; // input=-0.259765625, output=0.966450204846
			11'd1091: out = 32'b00000000000000000111101110010100; // input=-0.263671875, output=0.965439497855
			11'd1092: out = 32'b00000000000000000111101101110010; // input=-0.267578125, output=0.964414059445
			11'd1093: out = 32'b00000000000000000111101101010000; // input=-0.271484375, output=0.963373905264
			11'd1094: out = 32'b00000000000000000111101100101101; // input=-0.275390625, output=0.962319051181
			11'd1095: out = 32'b00000000000000000111101100001010; // input=-0.279296875, output=0.961249513295
			11'd1096: out = 32'b00000000000000000111101011100111; // input=-0.283203125, output=0.960165307923
			11'd1097: out = 32'b00000000000000000111101011000011; // input=-0.287109375, output=0.95906645161
			11'd1098: out = 32'b00000000000000000111101010011110; // input=-0.291015625, output=0.957952961123
			11'd1099: out = 32'b00000000000000000111101001111001; // input=-0.294921875, output=0.956824853452
			11'd1100: out = 32'b00000000000000000111101001010100; // input=-0.298828125, output=0.955682145811
			11'd1101: out = 32'b00000000000000000111101000101110; // input=-0.302734375, output=0.954524855637
			11'd1102: out = 32'b00000000000000000111101000000111; // input=-0.306640625, output=0.953353000587
			11'd1103: out = 32'b00000000000000000111100111100001; // input=-0.310546875, output=0.952166598544
			11'd1104: out = 32'b00000000000000000111100110111001; // input=-0.314453125, output=0.95096566761
			11'd1105: out = 32'b00000000000000000111100110010001; // input=-0.318359375, output=0.94975022611
			11'd1106: out = 32'b00000000000000000111100101101001; // input=-0.322265625, output=0.94852029259
			11'd1107: out = 32'b00000000000000000111100101000000; // input=-0.326171875, output=0.947275885817
			11'd1108: out = 32'b00000000000000000111100100010111; // input=-0.330078125, output=0.94601702478
			11'd1109: out = 32'b00000000000000000111100011101101; // input=-0.333984375, output=0.944743728687
			11'd1110: out = 32'b00000000000000000111100011000011; // input=-0.337890625, output=0.943456016966
			11'd1111: out = 32'b00000000000000000111100010011000; // input=-0.341796875, output=0.942153909268
			11'd1112: out = 32'b00000000000000000111100001101101; // input=-0.345703125, output=0.940837425461
			11'd1113: out = 32'b00000000000000000111100001000010; // input=-0.349609375, output=0.939506585632
			11'd1114: out = 32'b00000000000000000111100000010110; // input=-0.353515625, output=0.938161410088
			11'd1115: out = 32'b00000000000000000111011111101001; // input=-0.357421875, output=0.936801919355
			11'd1116: out = 32'b00000000000000000111011110111100; // input=-0.361328125, output=0.935428134178
			11'd1117: out = 32'b00000000000000000111011110001111; // input=-0.365234375, output=0.934040075518
			11'd1118: out = 32'b00000000000000000111011101100001; // input=-0.369140625, output=0.932637764556
			11'd1119: out = 32'b00000000000000000111011100110010; // input=-0.373046875, output=0.931221222689
			11'd1120: out = 32'b00000000000000000111011100000011; // input=-0.376953125, output=0.929790471532
			11'd1121: out = 32'b00000000000000000111011011010100; // input=-0.380859375, output=0.928345532916
			11'd1122: out = 32'b00000000000000000111011010100100; // input=-0.384765625, output=0.92688642889
			11'd1123: out = 32'b00000000000000000111011001110100; // input=-0.388671875, output=0.925413181717
			11'd1124: out = 32'b00000000000000000111011001000011; // input=-0.392578125, output=0.923925813877
			11'd1125: out = 32'b00000000000000000111011000010010; // input=-0.396484375, output=0.922424348067
			11'd1126: out = 32'b00000000000000000111010111100000; // input=-0.400390625, output=0.920908807195
			11'd1127: out = 32'b00000000000000000111010110101110; // input=-0.404296875, output=0.919379214389
			11'd1128: out = 32'b00000000000000000111010101111100; // input=-0.408203125, output=0.917835592986
			11'd1129: out = 32'b00000000000000000111010101001001; // input=-0.412109375, output=0.916277966542
			11'd1130: out = 32'b00000000000000000111010100010101; // input=-0.416015625, output=0.914706358823
			11'd1131: out = 32'b00000000000000000111010011100001; // input=-0.419921875, output=0.913120793811
			11'd1132: out = 32'b00000000000000000111010010101101; // input=-0.423828125, output=0.911521295699
			11'd1133: out = 32'b00000000000000000111010001111000; // input=-0.427734375, output=0.909907888893
			11'd1134: out = 32'b00000000000000000111010001000011; // input=-0.431640625, output=0.908280598013
			11'd1135: out = 32'b00000000000000000111010000001101; // input=-0.435546875, output=0.906639447888
			11'd1136: out = 32'b00000000000000000111001111010111; // input=-0.439453125, output=0.90498446356
			11'd1137: out = 32'b00000000000000000111001110100000; // input=-0.443359375, output=0.903315670283
			11'd1138: out = 32'b00000000000000000111001101101001; // input=-0.447265625, output=0.901633093521
			11'd1139: out = 32'b00000000000000000111001100110001; // input=-0.451171875, output=0.899936758946
			11'd1140: out = 32'b00000000000000000111001011111001; // input=-0.455078125, output=0.898226692444
			11'd1141: out = 32'b00000000000000000111001011000001; // input=-0.458984375, output=0.896502920108
			11'd1142: out = 32'b00000000000000000111001010001000; // input=-0.462890625, output=0.89476546824
			11'd1143: out = 32'b00000000000000000111001001001110; // input=-0.466796875, output=0.893014363352
			11'd1144: out = 32'b00000000000000000111001000010100; // input=-0.470703125, output=0.891249632163
			11'd1145: out = 32'b00000000000000000111000111011010; // input=-0.474609375, output=0.889471301602
			11'd1146: out = 32'b00000000000000000111000110011111; // input=-0.478515625, output=0.887679398803
			11'd1147: out = 32'b00000000000000000111000101100100; // input=-0.482421875, output=0.885873951108
			11'd1148: out = 32'b00000000000000000111000100101001; // input=-0.486328125, output=0.884054986067
			11'd1149: out = 32'b00000000000000000111000011101101; // input=-0.490234375, output=0.882222531435
			11'd1150: out = 32'b00000000000000000111000010110000; // input=-0.494140625, output=0.880376615172
			11'd1151: out = 32'b00000000000000000111000001110011; // input=-0.498046875, output=0.878517265445
			11'd1152: out = 32'b00000000000000000111000000110110; // input=-0.501953125, output=0.876644510625
			11'd1153: out = 32'b00000000000000000110111111111000; // input=-0.505859375, output=0.874758379289
			11'd1154: out = 32'b00000000000000000110111110111010; // input=-0.509765625, output=0.872858900216
			11'd1155: out = 32'b00000000000000000110111101111011; // input=-0.513671875, output=0.870946102391
			11'd1156: out = 32'b00000000000000000110111100111100; // input=-0.517578125, output=0.869020014999
			11'd1157: out = 32'b00000000000000000110111011111100; // input=-0.521484375, output=0.867080667431
			11'd1158: out = 32'b00000000000000000110111010111101; // input=-0.525390625, output=0.865128089279
			11'd1159: out = 32'b00000000000000000110111001111100; // input=-0.529296875, output=0.863162310337
			11'd1160: out = 32'b00000000000000000110111000111011; // input=-0.533203125, output=0.861183360599
			11'd1161: out = 32'b00000000000000000110110111111010; // input=-0.537109375, output=0.859191270264
			11'd1162: out = 32'b00000000000000000110110110111000; // input=-0.541015625, output=0.857186069726
			11'd1163: out = 32'b00000000000000000110110101110110; // input=-0.544921875, output=0.855167789584
			11'd1164: out = 32'b00000000000000000110110100110100; // input=-0.548828125, output=0.853136460634
			11'd1165: out = 32'b00000000000000000110110011110001; // input=-0.552734375, output=0.85109211387
			11'd1166: out = 32'b00000000000000000110110010101101; // input=-0.556640625, output=0.849034780489
			11'd1167: out = 32'b00000000000000000110110001101001; // input=-0.560546875, output=0.846964491881
			11'd1168: out = 32'b00000000000000000110110000100101; // input=-0.564453125, output=0.844881279637
			11'd1169: out = 32'b00000000000000000110101111100000; // input=-0.568359375, output=0.842785175544
			11'd1170: out = 32'b00000000000000000110101110011011; // input=-0.572265625, output=0.840676211586
			11'd1171: out = 32'b00000000000000000110101101010110; // input=-0.576171875, output=0.838554419944
			11'd1172: out = 32'b00000000000000000110101100010000; // input=-0.580078125, output=0.836419832992
			11'd1173: out = 32'b00000000000000000110101011001001; // input=-0.583984375, output=0.834272483304
			11'd1174: out = 32'b00000000000000000110101010000011; // input=-0.587890625, output=0.832112403643
			11'd1175: out = 32'b00000000000000000110101000111011; // input=-0.591796875, output=0.829939626972
			11'd1176: out = 32'b00000000000000000110100111110100; // input=-0.595703125, output=0.827754186442
			11'd1177: out = 32'b00000000000000000110100110101100; // input=-0.599609375, output=0.825556115402
			11'd1178: out = 32'b00000000000000000110100101100011; // input=-0.603515625, output=0.823345447392
			11'd1179: out = 32'b00000000000000000110100100011011; // input=-0.607421875, output=0.821122216143
			11'd1180: out = 32'b00000000000000000110100011010001; // input=-0.611328125, output=0.818886455579
			11'd1181: out = 32'b00000000000000000110100010001000; // input=-0.615234375, output=0.816638199815
			11'd1182: out = 32'b00000000000000000110100000111110; // input=-0.619140625, output=0.814377483157
			11'd1183: out = 32'b00000000000000000110011111110011; // input=-0.623046875, output=0.812104340101
			11'd1184: out = 32'b00000000000000000110011110101000; // input=-0.626953125, output=0.809818805332
			11'd1185: out = 32'b00000000000000000110011101011101; // input=-0.630859375, output=0.807520913724
			11'd1186: out = 32'b00000000000000000110011100010001; // input=-0.634765625, output=0.80521070034
			11'd1187: out = 32'b00000000000000000110011011000101; // input=-0.638671875, output=0.802888200432
			11'd1188: out = 32'b00000000000000000110011001111001; // input=-0.642578125, output=0.800553449438
			11'd1189: out = 32'b00000000000000000110011000101100; // input=-0.646484375, output=0.798206482983
			11'd1190: out = 32'b00000000000000000110010111011110; // input=-0.650390625, output=0.795847336879
			11'd1191: out = 32'b00000000000000000110010110010001; // input=-0.654296875, output=0.793476047124
			11'd1192: out = 32'b00000000000000000110010101000011; // input=-0.658203125, output=0.791092649901
			11'd1193: out = 32'b00000000000000000110010011110100; // input=-0.662109375, output=0.788697181577
			11'd1194: out = 32'b00000000000000000110010010100101; // input=-0.666015625, output=0.786289678704
			11'd1195: out = 32'b00000000000000000110010001010110; // input=-0.669921875, output=0.783870178019
			11'd1196: out = 32'b00000000000000000110010000000110; // input=-0.673828125, output=0.781438716439
			11'd1197: out = 32'b00000000000000000110001110110110; // input=-0.677734375, output=0.778995331066
			11'd1198: out = 32'b00000000000000000110001101100110; // input=-0.681640625, output=0.776540059182
			11'd1199: out = 32'b00000000000000000110001100010101; // input=-0.685546875, output=0.774072938252
			11'd1200: out = 32'b00000000000000000110001011000100; // input=-0.689453125, output=0.771594005922
			11'd1201: out = 32'b00000000000000000110001001110010; // input=-0.693359375, output=0.769103300017
			11'd1202: out = 32'b00000000000000000110001000100000; // input=-0.697265625, output=0.766600858541
			11'd1203: out = 32'b00000000000000000110000111001110; // input=-0.701171875, output=0.76408671968
			11'd1204: out = 32'b00000000000000000110000101111011; // input=-0.705078125, output=0.761560921795
			11'd1205: out = 32'b00000000000000000110000100101000; // input=-0.708984375, output=0.759023503428
			11'd1206: out = 32'b00000000000000000110000011010100; // input=-0.712890625, output=0.756474503295
			11'd1207: out = 32'b00000000000000000110000010000000; // input=-0.716796875, output=0.753913960293
			11'd1208: out = 32'b00000000000000000110000000101100; // input=-0.720703125, output=0.751341913491
			11'd1209: out = 32'b00000000000000000101111111010111; // input=-0.724609375, output=0.748758402136
			11'd1210: out = 32'b00000000000000000101111110000010; // input=-0.728515625, output=0.746163465649
			11'd1211: out = 32'b00000000000000000101111100101101; // input=-0.732421875, output=0.743557143625
			11'd1212: out = 32'b00000000000000000101111011010111; // input=-0.736328125, output=0.740939475835
			11'd1213: out = 32'b00000000000000000101111010000001; // input=-0.740234375, output=0.738310502219
			11'd1214: out = 32'b00000000000000000101111000101010; // input=-0.744140625, output=0.735670262894
			11'd1215: out = 32'b00000000000000000101110111010100; // input=-0.748046875, output=0.733018798145
			11'd1216: out = 32'b00000000000000000101110101111100; // input=-0.751953125, output=0.730356148432
			11'd1217: out = 32'b00000000000000000101110100100101; // input=-0.755859375, output=0.727682354382
			11'd1218: out = 32'b00000000000000000101110011001101; // input=-0.759765625, output=0.724997456795
			11'd1219: out = 32'b00000000000000000101110001110100; // input=-0.763671875, output=0.722301496639
			11'd1220: out = 32'b00000000000000000101110000011100; // input=-0.767578125, output=0.71959451505
			11'd1221: out = 32'b00000000000000000101101111000011; // input=-0.771484375, output=0.716876553335
			11'd1222: out = 32'b00000000000000000101101101101001; // input=-0.775390625, output=0.714147652965
			11'd1223: out = 32'b00000000000000000101101100001111; // input=-0.779296875, output=0.711407855581
			11'd1224: out = 32'b00000000000000000101101010110101; // input=-0.783203125, output=0.708657202988
			11'd1225: out = 32'b00000000000000000101101001011011; // input=-0.787109375, output=0.705895737158
			11'd1226: out = 32'b00000000000000000101101000000000; // input=-0.791015625, output=0.703123500228
			11'd1227: out = 32'b00000000000000000101100110100101; // input=-0.794921875, output=0.700340534498
			11'd1228: out = 32'b00000000000000000101100101001001; // input=-0.798828125, output=0.697546882433
			11'd1229: out = 32'b00000000000000000101100011101101; // input=-0.802734375, output=0.694742586661
			11'd1230: out = 32'b00000000000000000101100010010001; // input=-0.806640625, output=0.691927689972
			11'd1231: out = 32'b00000000000000000101100000110101; // input=-0.810546875, output=0.689102235318
			11'd1232: out = 32'b00000000000000000101011111011000; // input=-0.814453125, output=0.686266265812
			11'd1233: out = 32'b00000000000000000101011101111010; // input=-0.818359375, output=0.683419824726
			11'd1234: out = 32'b00000000000000000101011100011101; // input=-0.822265625, output=0.680562955495
			11'd1235: out = 32'b00000000000000000101011010111111; // input=-0.826171875, output=0.677695701711
			11'd1236: out = 32'b00000000000000000101011001100000; // input=-0.830078125, output=0.674818107123
			11'd1237: out = 32'b00000000000000000101011000000010; // input=-0.833984375, output=0.671930215642
			11'd1238: out = 32'b00000000000000000101010110100011; // input=-0.837890625, output=0.669032071333
			11'd1239: out = 32'b00000000000000000101010101000100; // input=-0.841796875, output=0.666123718417
			11'd1240: out = 32'b00000000000000000101010011100100; // input=-0.845703125, output=0.663205201273
			11'd1241: out = 32'b00000000000000000101010010000100; // input=-0.849609375, output=0.660276564433
			11'd1242: out = 32'b00000000000000000101010000100100; // input=-0.853515625, output=0.657337852585
			11'd1243: out = 32'b00000000000000000101001111000011; // input=-0.857421875, output=0.654389110571
			11'd1244: out = 32'b00000000000000000101001101100010; // input=-0.861328125, output=0.651430383384
			11'd1245: out = 32'b00000000000000000101001100000001; // input=-0.865234375, output=0.64846171617
			11'd1246: out = 32'b00000000000000000101001010011111; // input=-0.869140625, output=0.645483154229
			11'd1247: out = 32'b00000000000000000101001000111101; // input=-0.873046875, output=0.642494743009
			11'd1248: out = 32'b00000000000000000101000111011011; // input=-0.876953125, output=0.63949652811
			11'd1249: out = 32'b00000000000000000101000101111000; // input=-0.880859375, output=0.63648855528
			11'd1250: out = 32'b00000000000000000101000100010110; // input=-0.884765625, output=0.633470870418
			11'd1251: out = 32'b00000000000000000101000010110010; // input=-0.888671875, output=0.63044351957
			11'd1252: out = 32'b00000000000000000101000001001111; // input=-0.892578125, output=0.62740654893
			11'd1253: out = 32'b00000000000000000100111111101011; // input=-0.896484375, output=0.624360004837
			11'd1254: out = 32'b00000000000000000100111110000111; // input=-0.900390625, output=0.621303933779
			11'd1255: out = 32'b00000000000000000100111100100010; // input=-0.904296875, output=0.618238382388
			11'd1256: out = 32'b00000000000000000100111010111110; // input=-0.908203125, output=0.615163397439
			11'd1257: out = 32'b00000000000000000100111001011001; // input=-0.912109375, output=0.612079025854
			11'd1258: out = 32'b00000000000000000100110111110011; // input=-0.916015625, output=0.608985314696
			11'd1259: out = 32'b00000000000000000100110110001110; // input=-0.919921875, output=0.605882311171
			11'd1260: out = 32'b00000000000000000100110100101000; // input=-0.923828125, output=0.602770062628
			11'd1261: out = 32'b00000000000000000100110011000001; // input=-0.927734375, output=0.599648616555
			11'd1262: out = 32'b00000000000000000100110001011011; // input=-0.931640625, output=0.596518020582
			11'd1263: out = 32'b00000000000000000100101111110100; // input=-0.935546875, output=0.593378322478
			11'd1264: out = 32'b00000000000000000100101110001101; // input=-0.939453125, output=0.590229570151
			11'd1265: out = 32'b00000000000000000100101100100101; // input=-0.943359375, output=0.587071811646
			11'd1266: out = 32'b00000000000000000100101010111101; // input=-0.947265625, output=0.583905095149
			11'd1267: out = 32'b00000000000000000100101001010101; // input=-0.951171875, output=0.580729468977
			11'd1268: out = 32'b00000000000000000100100111101101; // input=-0.955078125, output=0.577544981589
			11'd1269: out = 32'b00000000000000000100100110000100; // input=-0.958984375, output=0.574351681575
			11'd1270: out = 32'b00000000000000000100100100011011; // input=-0.962890625, output=0.571149617661
			11'd1271: out = 32'b00000000000000000100100010110010; // input=-0.966796875, output=0.567938838706
			11'd1272: out = 32'b00000000000000000100100001001001; // input=-0.970703125, output=0.564719393703
			11'd1273: out = 32'b00000000000000000100011111011111; // input=-0.974609375, output=0.561491331777
			11'd1274: out = 32'b00000000000000000100011101110101; // input=-0.978515625, output=0.558254702185
			11'd1275: out = 32'b00000000000000000100011100001011; // input=-0.982421875, output=0.555009554312
			11'd1276: out = 32'b00000000000000000100011010100000; // input=-0.986328125, output=0.551755937677
			11'd1277: out = 32'b00000000000000000100011000110101; // input=-0.990234375, output=0.548493901924
			11'd1278: out = 32'b00000000000000000100010111001010; // input=-0.994140625, output=0.54522349683
			11'd1279: out = 32'b00000000000000000100010101011110; // input=-0.998046875, output=0.541944772296
			11'd1280: out = 32'b00000000000000000100010011110011; // input=-1.001953125, output=0.538657778351
			11'd1281: out = 32'b00000000000000000100010010000111; // input=-1.005859375, output=0.535362565152
			11'd1282: out = 32'b00000000000000000100010000011011; // input=-1.009765625, output=0.532059182978
			11'd1283: out = 32'b00000000000000000100001110101110; // input=-1.013671875, output=0.528747682236
			11'd1284: out = 32'b00000000000000000100001101000001; // input=-1.017578125, output=0.525428113455
			11'd1285: out = 32'b00000000000000000100001011010100; // input=-1.021484375, output=0.522100527287
			11'd1286: out = 32'b00000000000000000100001001100111; // input=-1.025390625, output=0.518764974507
			11'd1287: out = 32'b00000000000000000100000111111001; // input=-1.029296875, output=0.515421506013
			11'd1288: out = 32'b00000000000000000100000110001100; // input=-1.033203125, output=0.51207017282
			11'd1289: out = 32'b00000000000000000100000100011101; // input=-1.037109375, output=0.508711026066
			11'd1290: out = 32'b00000000000000000100000010101111; // input=-1.041015625, output=0.505344117008
			11'd1291: out = 32'b00000000000000000100000001000001; // input=-1.044921875, output=0.501969497021
			11'd1292: out = 32'b00000000000000000011111111010010; // input=-1.048828125, output=0.498587217597
			11'd1293: out = 32'b00000000000000000011111101100011; // input=-1.052734375, output=0.495197330345
			11'd1294: out = 32'b00000000000000000011111011110011; // input=-1.056640625, output=0.491799886991
			11'd1295: out = 32'b00000000000000000011111010000100; // input=-1.060546875, output=0.488394939376
			11'd1296: out = 32'b00000000000000000011111000010100; // input=-1.064453125, output=0.484982539455
			11'd1297: out = 32'b00000000000000000011110110100100; // input=-1.068359375, output=0.481562739297
			11'd1298: out = 32'b00000000000000000011110100110100; // input=-1.072265625, output=0.478135591084
			11'd1299: out = 32'b00000000000000000011110011000011; // input=-1.076171875, output=0.474701147111
			11'd1300: out = 32'b00000000000000000011110001010010; // input=-1.080078125, output=0.471259459782
			11'd1301: out = 32'b00000000000000000011101111100001; // input=-1.083984375, output=0.467810581613
			11'd1302: out = 32'b00000000000000000011101101110000; // input=-1.087890625, output=0.464354565231
			11'd1303: out = 32'b00000000000000000011101011111110; // input=-1.091796875, output=0.460891463369
			11'd1304: out = 32'b00000000000000000011101010001101; // input=-1.095703125, output=0.45742132887
			11'd1305: out = 32'b00000000000000000011101000011011; // input=-1.099609375, output=0.453944214685
			11'd1306: out = 32'b00000000000000000011100110101001; // input=-1.103515625, output=0.45046017387
			11'd1307: out = 32'b00000000000000000011100100110110; // input=-1.107421875, output=0.446969259586
			11'd1308: out = 32'b00000000000000000011100011000100; // input=-1.111328125, output=0.443471525102
			11'd1309: out = 32'b00000000000000000011100001010001; // input=-1.115234375, output=0.439967023787
			11'd1310: out = 32'b00000000000000000011011111011110; // input=-1.119140625, output=0.436455809118
			11'd1311: out = 32'b00000000000000000011011101101011; // input=-1.123046875, output=0.432937934669
			11'd1312: out = 32'b00000000000000000011011011110111; // input=-1.126953125, output=0.429413454121
			11'd1313: out = 32'b00000000000000000011011010000011; // input=-1.130859375, output=0.425882421251
			11'd1314: out = 32'b00000000000000000011011000001111; // input=-1.134765625, output=0.42234488994
			11'd1315: out = 32'b00000000000000000011010110011011; // input=-1.138671875, output=0.418800914165
			11'd1316: out = 32'b00000000000000000011010100100111; // input=-1.142578125, output=0.415250548003
			11'd1317: out = 32'b00000000000000000011010010110010; // input=-1.146484375, output=0.411693845629
			11'd1318: out = 32'b00000000000000000011010000111110; // input=-1.150390625, output=0.408130861314
			11'd1319: out = 32'b00000000000000000011001111001001; // input=-1.154296875, output=0.404561649424
			11'd1320: out = 32'b00000000000000000011001101010100; // input=-1.158203125, output=0.40098626442
			11'd1321: out = 32'b00000000000000000011001011011110; // input=-1.162109375, output=0.39740476086
			11'd1322: out = 32'b00000000000000000011001001101001; // input=-1.166015625, output=0.393817193392
			11'd1323: out = 32'b00000000000000000011000111110011; // input=-1.169921875, output=0.390223616758
			11'd1324: out = 32'b00000000000000000011000101111101; // input=-1.173828125, output=0.386624085792
			11'd1325: out = 32'b00000000000000000011000100000111; // input=-1.177734375, output=0.383018655418
			11'd1326: out = 32'b00000000000000000011000010010000; // input=-1.181640625, output=0.37940738065
			11'd1327: out = 32'b00000000000000000011000000011010; // input=-1.185546875, output=0.375790316593
			11'd1328: out = 32'b00000000000000000010111110100011; // input=-1.189453125, output=0.372167518438
			11'd1329: out = 32'b00000000000000000010111100101100; // input=-1.193359375, output=0.368539041464
			11'd1330: out = 32'b00000000000000000010111010110101; // input=-1.197265625, output=0.364904941038
			11'd1331: out = 32'b00000000000000000010111000111110; // input=-1.201171875, output=0.361265272612
			11'd1332: out = 32'b00000000000000000010110111000110; // input=-1.205078125, output=0.357620091721
			11'd1333: out = 32'b00000000000000000010110101001111; // input=-1.208984375, output=0.353969453989
			11'd1334: out = 32'b00000000000000000010110011010111; // input=-1.212890625, output=0.350313415118
			11'd1335: out = 32'b00000000000000000010110001011111; // input=-1.216796875, output=0.346652030895
			11'd1336: out = 32'b00000000000000000010101111100111; // input=-1.220703125, output=0.342985357189
			11'd1337: out = 32'b00000000000000000010101101101111; // input=-1.224609375, output=0.339313449948
			11'd1338: out = 32'b00000000000000000010101011110110; // input=-1.228515625, output=0.335636365202
			11'd1339: out = 32'b00000000000000000010101001111101; // input=-1.232421875, output=0.331954159057
			11'd1340: out = 32'b00000000000000000010101000000101; // input=-1.236328125, output=0.328266887701
			11'd1341: out = 32'b00000000000000000010100110001100; // input=-1.240234375, output=0.324574607395
			11'd1342: out = 32'b00000000000000000010100100010011; // input=-1.244140625, output=0.320877374481
			11'd1343: out = 32'b00000000000000000010100010011001; // input=-1.248046875, output=0.317175245372
			11'd1344: out = 32'b00000000000000000010100000100000; // input=-1.251953125, output=0.31346827656
			11'd1345: out = 32'b00000000000000000010011110100110; // input=-1.255859375, output=0.309756524607
			11'd1346: out = 32'b00000000000000000010011100101100; // input=-1.259765625, output=0.306040046151
			11'd1347: out = 32'b00000000000000000010011010110010; // input=-1.263671875, output=0.3023188979
			11'd1348: out = 32'b00000000000000000010011000111000; // input=-1.267578125, output=0.298593136635
			11'd1349: out = 32'b00000000000000000010010110111110; // input=-1.271484375, output=0.294862819205
			11'd1350: out = 32'b00000000000000000010010101000100; // input=-1.275390625, output=0.291128002532
			11'd1351: out = 32'b00000000000000000010010011001001; // input=-1.279296875, output=0.287388743604
			11'd1352: out = 32'b00000000000000000010010001001110; // input=-1.283203125, output=0.283645099478
			11'd1353: out = 32'b00000000000000000010001111010100; // input=-1.287109375, output=0.279897127276
			11'd1354: out = 32'b00000000000000000010001101011001; // input=-1.291015625, output=0.276144884188
			11'd1355: out = 32'b00000000000000000010001011011110; // input=-1.294921875, output=0.272388427469
			11'd1356: out = 32'b00000000000000000010001001100010; // input=-1.298828125, output=0.268627814438
			11'd1357: out = 32'b00000000000000000010000111100111; // input=-1.302734375, output=0.264863102477
			11'd1358: out = 32'b00000000000000000010000101101100; // input=-1.306640625, output=0.26109434903
			11'd1359: out = 32'b00000000000000000010000011110000; // input=-1.310546875, output=0.257321611606
			11'd1360: out = 32'b00000000000000000010000001110100; // input=-1.314453125, output=0.25354494777
			11'd1361: out = 32'b00000000000000000001111111111000; // input=-1.318359375, output=0.24976441515
			11'd1362: out = 32'b00000000000000000001111101111100; // input=-1.322265625, output=0.245980071432
			11'd1363: out = 32'b00000000000000000001111100000000; // input=-1.326171875, output=0.242191974361
			11'd1364: out = 32'b00000000000000000001111010000100; // input=-1.330078125, output=0.238400181739
			11'd1365: out = 32'b00000000000000000001111000001000; // input=-1.333984375, output=0.234604751423
			11'd1366: out = 32'b00000000000000000001110110001011; // input=-1.337890625, output=0.230805741327
			11'd1367: out = 32'b00000000000000000001110100001110; // input=-1.341796875, output=0.22700320942
			11'd1368: out = 32'b00000000000000000001110010010010; // input=-1.345703125, output=0.223197213723
			11'd1369: out = 32'b00000000000000000001110000010101; // input=-1.349609375, output=0.219387812311
			11'd1370: out = 32'b00000000000000000001101110011000; // input=-1.353515625, output=0.215575063311
			11'd1371: out = 32'b00000000000000000001101100011011; // input=-1.357421875, output=0.211759024901
			11'd1372: out = 32'b00000000000000000001101010011110; // input=-1.361328125, output=0.207939755308
			11'd1373: out = 32'b00000000000000000001101000100001; // input=-1.365234375, output=0.204117312811
			11'd1374: out = 32'b00000000000000000001100110100011; // input=-1.369140625, output=0.200291755735
			11'd1375: out = 32'b00000000000000000001100100100110; // input=-1.373046875, output=0.196463142453
			11'd1376: out = 32'b00000000000000000001100010101000; // input=-1.376953125, output=0.192631531385
			11'd1377: out = 32'b00000000000000000001100000101010; // input=-1.380859375, output=0.188796980997
			11'd1378: out = 32'b00000000000000000001011110101101; // input=-1.384765625, output=0.184959549799
			11'd1379: out = 32'b00000000000000000001011100101111; // input=-1.388671875, output=0.181119296346
			11'd1380: out = 32'b00000000000000000001011010110001; // input=-1.392578125, output=0.177276279236
			11'd1381: out = 32'b00000000000000000001011000110011; // input=-1.396484375, output=0.173430557107
			11'd1382: out = 32'b00000000000000000001010110110101; // input=-1.400390625, output=0.169582188642
			11'd1383: out = 32'b00000000000000000001010100110111; // input=-1.404296875, output=0.165731232561
			11'd1384: out = 32'b00000000000000000001010010111000; // input=-1.408203125, output=0.161877747625
			11'd1385: out = 32'b00000000000000000001010000111010; // input=-1.412109375, output=0.158021792634
			11'd1386: out = 32'b00000000000000000001001110111100; // input=-1.416015625, output=0.154163426425
			11'd1387: out = 32'b00000000000000000001001100111101; // input=-1.419921875, output=0.150302707872
			11'd1388: out = 32'b00000000000000000001001010111111; // input=-1.423828125, output=0.146439695884
			11'd1389: out = 32'b00000000000000000001001001000000; // input=-1.427734375, output=0.142574449407
			11'd1390: out = 32'b00000000000000000001000111000001; // input=-1.431640625, output=0.138707027419
			11'd1391: out = 32'b00000000000000000001000101000010; // input=-1.435546875, output=0.134837488933
			11'd1392: out = 32'b00000000000000000001000011000011; // input=-1.439453125, output=0.130965892992
			11'd1393: out = 32'b00000000000000000001000001000101; // input=-1.443359375, output=0.127092298673
			11'd1394: out = 32'b00000000000000000000111111000110; // input=-1.447265625, output=0.123216765082
			11'd1395: out = 32'b00000000000000000000111101000111; // input=-1.451171875, output=0.119339351355
			11'd1396: out = 32'b00000000000000000000111011000111; // input=-1.455078125, output=0.115460116656
			11'd1397: out = 32'b00000000000000000000111001001000; // input=-1.458984375, output=0.111579120177
			11'd1398: out = 32'b00000000000000000000110111001001; // input=-1.462890625, output=0.107696421139
			11'd1399: out = 32'b00000000000000000000110101001010; // input=-1.466796875, output=0.103812078785
			11'd1400: out = 32'b00000000000000000000110011001010; // input=-1.470703125, output=0.0999261523872
			11'd1401: out = 32'b00000000000000000000110001001011; // input=-1.474609375, output=0.0960387012391
			11'd1402: out = 32'b00000000000000000000101111001100; // input=-1.478515625, output=0.0921497846586
			11'd1403: out = 32'b00000000000000000000101101001100; // input=-1.482421875, output=0.0882594619857
			11'd1404: out = 32'b00000000000000000000101011001101; // input=-1.486328125, output=0.084367792582
			11'd1405: out = 32'b00000000000000000000101001001101; // input=-1.490234375, output=0.0804748358296
			11'd1406: out = 32'b00000000000000000000100111001101; // input=-1.494140625, output=0.0765806511302
			11'd1407: out = 32'b00000000000000000000100101001110; // input=-1.498046875, output=0.0726852979043
			11'd1408: out = 32'b00000000000000000000100011001110; // input=-1.501953125, output=0.0687888355902
			11'd1409: out = 32'b00000000000000000000100001001110; // input=-1.505859375, output=0.0648913236431
			11'd1410: out = 32'b00000000000000000000011111001111; // input=-1.509765625, output=0.0609928215342
			11'd1411: out = 32'b00000000000000000000011101001111; // input=-1.513671875, output=0.0570933887499
			11'd1412: out = 32'b00000000000000000000011011001111; // input=-1.517578125, output=0.0531930847907
			11'd1413: out = 32'b00000000000000000000011001001111; // input=-1.521484375, output=0.0492919691706
			11'd1414: out = 32'b00000000000000000000010111001111; // input=-1.525390625, output=0.0453901014156
			11'd1415: out = 32'b00000000000000000000010101001111; // input=-1.529296875, output=0.0414875410635
			11'd1416: out = 32'b00000000000000000000010011010000; // input=-1.533203125, output=0.0375843476626
			11'd1417: out = 32'b00000000000000000000010001010000; // input=-1.537109375, output=0.0336805807707
			11'd1418: out = 32'b00000000000000000000001111010000; // input=-1.541015625, output=0.0297762999547
			11'd1419: out = 32'b00000000000000000000001101010000; // input=-1.544921875, output=0.0258715647889
			11'd1420: out = 32'b00000000000000000000001011010000; // input=-1.548828125, output=0.0219664348549
			11'd1421: out = 32'b00000000000000000000001001010000; // input=-1.552734375, output=0.0180609697401
			11'd1422: out = 32'b00000000000000000000000111010000; // input=-1.556640625, output=0.0141552290372
			11'd1423: out = 32'b00000000000000000000000101010000; // input=-1.560546875, output=0.0102492723429
			11'd1424: out = 32'b00000000000000000000000011010000; // input=-1.564453125, output=0.00634315925725
			11'd1425: out = 32'b00000000000000000000000001010000; // input=-1.568359375, output=0.00243694938283
			11'd1426: out = 32'b10000000000000000000000000110000; // input=-1.572265625, output=-0.00146929767644
			11'd1427: out = 32'b10000000000000000000000010110000; // input=-1.576171875, output=-0.00537552231604
			11'd1428: out = 32'b10000000000000000000000100110000; // input=-1.580078125, output=-0.00928166493177
			11'd1429: out = 32'b10000000000000000000000110110000; // input=-1.583984375, output=-0.0131876659207
			11'd1430: out = 32'b10000000000000000000001000110000; // input=-1.587890625, output=-0.0170934656821
			11'd1431: out = 32'b10000000000000000000001010110000; // input=-1.591796875, output=-0.0209990046183
			11'd1432: out = 32'b10000000000000000000001100110000; // input=-1.595703125, output=-0.0249042231354
			11'd1433: out = 32'b10000000000000000000001110110000; // input=-1.599609375, output=-0.0288090616448
			11'd1434: out = 32'b10000000000000000000010000110000; // input=-1.603515625, output=-0.0327134605633
			11'd1435: out = 32'b10000000000000000000010010110000; // input=-1.607421875, output=-0.0366173603147
			11'd1436: out = 32'b10000000000000000000010100110000; // input=-1.611328125, output=-0.0405207013302
			11'd1437: out = 32'b10000000000000000000010110110000; // input=-1.615234375, output=-0.0444234240496
			11'd1438: out = 32'b10000000000000000000011000110000; // input=-1.619140625, output=-0.0483254689223
			11'd1439: out = 32'b10000000000000000000011010101111; // input=-1.623046875, output=-0.0522267764077
			11'd1440: out = 32'b10000000000000000000011100101111; // input=-1.626953125, output=-0.0561272869768
			11'd1441: out = 32'b10000000000000000000011110101111; // input=-1.630859375, output=-0.0600269411126
			11'd1442: out = 32'b10000000000000000000100000101111; // input=-1.634765625, output=-0.0639256793111
			11'd1443: out = 32'b10000000000000000000100010101110; // input=-1.638671875, output=-0.0678234420824
			11'd1444: out = 32'b10000000000000000000100100101110; // input=-1.642578125, output=-0.0717201699514
			11'd1445: out = 32'b10000000000000000000100110101110; // input=-1.646484375, output=-0.0756158034588
			11'd1446: out = 32'b10000000000000000000101000101101; // input=-1.650390625, output=-0.0795102831621
			11'd1447: out = 32'b10000000000000000000101010101101; // input=-1.654296875, output=-0.0834035496363
			11'd1448: out = 32'b10000000000000000000101100101101; // input=-1.658203125, output=-0.087295543475
			11'd1449: out = 32'b10000000000000000000101110101100; // input=-1.662109375, output=-0.0911862052911
			11'd1450: out = 32'b10000000000000000000110000101011; // input=-1.666015625, output=-0.0950754757179
			11'd1451: out = 32'b10000000000000000000110010101011; // input=-1.669921875, output=-0.0989632954099
			11'd1452: out = 32'b10000000000000000000110100101010; // input=-1.673828125, output=-0.102849605044
			11'd1453: out = 32'b10000000000000000000110110101001; // input=-1.677734375, output=-0.106734345319
			11'd1454: out = 32'b10000000000000000000111000101001; // input=-1.681640625, output=-0.11061745696
			11'd1455: out = 32'b10000000000000000000111010101000; // input=-1.685546875, output=-0.114498880714
			11'd1456: out = 32'b10000000000000000000111100100111; // input=-1.689453125, output=-0.118378557356
			11'd1457: out = 32'b10000000000000000000111110100110; // input=-1.693359375, output=-0.122256427688
			11'd1458: out = 32'b10000000000000000001000000100101; // input=-1.697265625, output=-0.126132432536
			11'd1459: out = 32'b10000000000000000001000010100100; // input=-1.701171875, output=-0.130006512759
			11'd1460: out = 32'b10000000000000000001000100100011; // input=-1.705078125, output=-0.133878609242
			11'd1461: out = 32'b10000000000000000001000110100010; // input=-1.708984375, output=-0.137748662903
			11'd1462: out = 32'b10000000000000000001001000100000; // input=-1.712890625, output=-0.141616614688
			11'd1463: out = 32'b10000000000000000001001010011111; // input=-1.716796875, output=-0.145482405578
			11'd1464: out = 32'b10000000000000000001001100011110; // input=-1.720703125, output=-0.149345976585
			11'd1465: out = 32'b10000000000000000001001110011100; // input=-1.724609375, output=-0.153207268757
			11'd1466: out = 32'b10000000000000000001010000011011; // input=-1.728515625, output=-0.157066223174
			11'd1467: out = 32'b10000000000000000001010010011001; // input=-1.732421875, output=-0.160922780954
			11'd1468: out = 32'b10000000000000000001010100010111; // input=-1.736328125, output=-0.164776883251
			11'd1469: out = 32'b10000000000000000001010110010110; // input=-1.740234375, output=-0.168628471254
			11'd1470: out = 32'b10000000000000000001011000010100; // input=-1.744140625, output=-0.172477486195
			11'd1471: out = 32'b10000000000000000001011010010010; // input=-1.748046875, output=-0.176323869342
			11'd1472: out = 32'b10000000000000000001011100010000; // input=-1.751953125, output=-0.180167562003
			11'd1473: out = 32'b10000000000000000001011110001110; // input=-1.755859375, output=-0.184008505529
			11'd1474: out = 32'b10000000000000000001100000001011; // input=-1.759765625, output=-0.187846641311
			11'd1475: out = 32'b10000000000000000001100010001001; // input=-1.763671875, output=-0.191681910785
			11'd1476: out = 32'b10000000000000000001100100000111; // input=-1.767578125, output=-0.195514255429
			11'd1477: out = 32'b10000000000000000001100110000100; // input=-1.771484375, output=-0.199343616766
			11'd1478: out = 32'b10000000000000000001101000000001; // input=-1.775390625, output=-0.203169936364
			11'd1479: out = 32'b10000000000000000001101001111111; // input=-1.779296875, output=-0.206993155839
			11'd1480: out = 32'b10000000000000000001101011111100; // input=-1.783203125, output=-0.210813216853
			11'd1481: out = 32'b10000000000000000001101101111001; // input=-1.787109375, output=-0.214630061117
			11'd1482: out = 32'b10000000000000000001101111110110; // input=-1.791015625, output=-0.218443630391
			11'd1483: out = 32'b10000000000000000001110001110011; // input=-1.794921875, output=-0.222253866483
			11'd1484: out = 32'b10000000000000000001110011110000; // input=-1.798828125, output=-0.226060711255
			11'd1485: out = 32'b10000000000000000001110101101100; // input=-1.802734375, output=-0.229864106618
			11'd1486: out = 32'b10000000000000000001110111101001; // input=-1.806640625, output=-0.233663994538
			11'd1487: out = 32'b10000000000000000001111001100101; // input=-1.810546875, output=-0.237460317033
			11'd1488: out = 32'b10000000000000000001111011100001; // input=-1.814453125, output=-0.241253016175
			11'd1489: out = 32'b10000000000000000001111101011110; // input=-1.818359375, output=-0.245042034094
			11'd1490: out = 32'b10000000000000000001111111011010; // input=-1.822265625, output=-0.248827312972
			11'd1491: out = 32'b10000000000000000010000001010101; // input=-1.826171875, output=-0.252608795052
			11'd1492: out = 32'b10000000000000000010000011010001; // input=-1.830078125, output=-0.256386422632
			11'd1493: out = 32'b10000000000000000010000101001101; // input=-1.833984375, output=-0.260160138071
			11'd1494: out = 32'b10000000000000000010000111001000; // input=-1.837890625, output=-0.263929883786
			11'd1495: out = 32'b10000000000000000010001001000100; // input=-1.841796875, output=-0.267695602256
			11'd1496: out = 32'b10000000000000000010001010111111; // input=-1.845703125, output=-0.271457236021
			11'd1497: out = 32'b10000000000000000010001100111010; // input=-1.849609375, output=-0.275214727682
			11'd1498: out = 32'b10000000000000000010001110110101; // input=-1.853515625, output=-0.278968019905
			11'd1499: out = 32'b10000000000000000010010000110000; // input=-1.857421875, output=-0.282717055419
			11'd1500: out = 32'b10000000000000000010010010101011; // input=-1.861328125, output=-0.286461777019
			11'd1501: out = 32'b10000000000000000010010100100101; // input=-1.865234375, output=-0.290202127564
			11'd1502: out = 32'b10000000000000000010010110100000; // input=-1.869140625, output=-0.293938049982
			11'd1503: out = 32'b10000000000000000010011000011010; // input=-1.873046875, output=-0.297669487267
			11'd1504: out = 32'b10000000000000000010011010010100; // input=-1.876953125, output=-0.301396382482
			11'd1505: out = 32'b10000000000000000010011100001110; // input=-1.880859375, output=-0.305118678759
			11'd1506: out = 32'b10000000000000000010011110001000; // input=-1.884765625, output=-0.308836319301
			11'd1507: out = 32'b10000000000000000010100000000010; // input=-1.888671875, output=-0.31254924738
			11'd1508: out = 32'b10000000000000000010100001111011; // input=-1.892578125, output=-0.316257406342
			11'd1509: out = 32'b10000000000000000010100011110100; // input=-1.896484375, output=-0.319960739605
			11'd1510: out = 32'b10000000000000000010100101101110; // input=-1.900390625, output=-0.323659190661
			11'd1511: out = 32'b10000000000000000010100111100111; // input=-1.904296875, output=-0.327352703076
			11'd1512: out = 32'b10000000000000000010101001100000; // input=-1.908203125, output=-0.331041220491
			11'd1513: out = 32'b10000000000000000010101011011000; // input=-1.912109375, output=-0.334724686625
			11'd1514: out = 32'b10000000000000000010101101010001; // input=-1.916015625, output=-0.338403045272
			11'd1515: out = 32'b10000000000000000010101111001001; // input=-1.919921875, output=-0.342076240304
			11'd1516: out = 32'b10000000000000000010110001000001; // input=-1.923828125, output=-0.345744215674
			11'd1517: out = 32'b10000000000000000010110010111001; // input=-1.927734375, output=-0.349406915413
			11'd1518: out = 32'b10000000000000000010110100110001; // input=-1.931640625, output=-0.353064283632
			11'd1519: out = 32'b10000000000000000010110110101001; // input=-1.935546875, output=-0.356716264525
			11'd1520: out = 32'b10000000000000000010111000100000; // input=-1.939453125, output=-0.360362802366
			11'd1521: out = 32'b10000000000000000010111010011000; // input=-1.943359375, output=-0.364003841514
			11'd1522: out = 32'b10000000000000000010111100001111; // input=-1.947265625, output=-0.367639326412
			11'd1523: out = 32'b10000000000000000010111110000110; // input=-1.951171875, output=-0.371269201585
			11'd1524: out = 32'b10000000000000000010111111111101; // input=-1.955078125, output=-0.374893411648
			11'd1525: out = 32'b10000000000000000011000001110011; // input=-1.958984375, output=-0.378511901298
			11'd1526: out = 32'b10000000000000000011000011101001; // input=-1.962890625, output=-0.382124615322
			11'd1527: out = 32'b10000000000000000011000101100000; // input=-1.966796875, output=-0.385731498595
			11'd1528: out = 32'b10000000000000000011000111010110; // input=-1.970703125, output=-0.38933249608
			11'd1529: out = 32'b10000000000000000011001001001011; // input=-1.974609375, output=-0.392927552829
			11'd1530: out = 32'b10000000000000000011001011000001; // input=-1.978515625, output=-0.396516613988
			11'd1531: out = 32'b10000000000000000011001100110110; // input=-1.982421875, output=-0.400099624791
			11'd1532: out = 32'b10000000000000000011001110101100; // input=-1.986328125, output=-0.403676530566
			11'd1533: out = 32'b10000000000000000011010000100001; // input=-1.990234375, output=-0.407247276734
			11'd1534: out = 32'b10000000000000000011010010010101; // input=-1.994140625, output=-0.41081180881
			11'd1535: out = 32'b10000000000000000011010100001010; // input=-1.998046875, output=-0.414370072403
			11'd1536: out = 32'b10000000000000000011010101111110; // input=-2.001953125, output=-0.417922013218
			11'd1537: out = 32'b10000000000000000011010111110011; // input=-2.005859375, output=-0.421467577057
			11'd1538: out = 32'b10000000000000000011011001100111; // input=-2.009765625, output=-0.42500670982
			11'd1539: out = 32'b10000000000000000011011011011010; // input=-2.013671875, output=-0.428539357504
			11'd1540: out = 32'b10000000000000000011011101001110; // input=-2.017578125, output=-0.432065466204
			11'd1541: out = 32'b10000000000000000011011111000001; // input=-2.021484375, output=-0.435584982116
			11'd1542: out = 32'b10000000000000000011100000110100; // input=-2.025390625, output=-0.439097851538
			11'd1543: out = 32'b10000000000000000011100010100111; // input=-2.029296875, output=-0.442604020867
			11'd1544: out = 32'b10000000000000000011100100011010; // input=-2.033203125, output=-0.446103436603
			11'd1545: out = 32'b10000000000000000011100110001100; // input=-2.037109375, output=-0.449596045349
			11'd1546: out = 32'b10000000000000000011100111111111; // input=-2.041015625, output=-0.453081793813
			11'd1547: out = 32'b10000000000000000011101001110001; // input=-2.044921875, output=-0.456560628806
			11'd1548: out = 32'b10000000000000000011101011100010; // input=-2.048828125, output=-0.460032497246
			11'd1549: out = 32'b10000000000000000011101101010100; // input=-2.052734375, output=-0.463497346155
			11'd1550: out = 32'b10000000000000000011101111000101; // input=-2.056640625, output=-0.466955122666
			11'd1551: out = 32'b10000000000000000011110000110110; // input=-2.060546875, output=-0.470405774016
			11'd1552: out = 32'b10000000000000000011110010100111; // input=-2.064453125, output=-0.473849247552
			11'd1553: out = 32'b10000000000000000011110100011000; // input=-2.068359375, output=-0.477285490732
			11'd1554: out = 32'b10000000000000000011110110001000; // input=-2.072265625, output=-0.480714451123
			11'd1555: out = 32'b10000000000000000011110111111000; // input=-2.076171875, output=-0.484136076402
			11'd1556: out = 32'b10000000000000000011111001101000; // input=-2.080078125, output=-0.487550314361
			11'd1557: out = 32'b10000000000000000011111011011000; // input=-2.083984375, output=-0.490957112901
			11'd1558: out = 32'b10000000000000000011111101000111; // input=-2.087890625, output=-0.49435642004
			11'd1559: out = 32'b10000000000000000011111110110110; // input=-2.091796875, output=-0.497748183909
			11'd1560: out = 32'b10000000000000000100000000100101; // input=-2.095703125, output=-0.501132352752
			11'd1561: out = 32'b10000000000000000100000010010100; // input=-2.099609375, output=-0.504508874933
			11'd1562: out = 32'b10000000000000000100000100000010; // input=-2.103515625, output=-0.507877698929
			11'd1563: out = 32'b10000000000000000100000101110000; // input=-2.107421875, output=-0.511238773335
			11'd1564: out = 32'b10000000000000000100000111011110; // input=-2.111328125, output=-0.514592046868
			11'd1565: out = 32'b10000000000000000100001001001100; // input=-2.115234375, output=-0.517937468358
			11'd1566: out = 32'b10000000000000000100001010111001; // input=-2.119140625, output=-0.52127498676
			11'd1567: out = 32'b10000000000000000100001100100110; // input=-2.123046875, output=-0.524604551148
			11'd1568: out = 32'b10000000000000000100001110010011; // input=-2.126953125, output=-0.527926110715
			11'd1569: out = 32'b10000000000000000100010000000000; // input=-2.130859375, output=-0.531239614779
			11'd1570: out = 32'b10000000000000000100010001101100; // input=-2.134765625, output=-0.53454501278
			11'd1571: out = 32'b10000000000000000100010011011000; // input=-2.138671875, output=-0.537842254283
			11'd1572: out = 32'b10000000000000000100010101000100; // input=-2.142578125, output=-0.541131288974
			11'd1573: out = 32'b10000000000000000100010110101111; // input=-2.146484375, output=-0.544412066667
			11'd1574: out = 32'b10000000000000000100011000011011; // input=-2.150390625, output=-0.547684537302
			11'd1575: out = 32'b10000000000000000100011010000101; // input=-2.154296875, output=-0.550948650945
			11'd1576: out = 32'b10000000000000000100011011110000; // input=-2.158203125, output=-0.554204357789
			11'd1577: out = 32'b10000000000000000100011101011011; // input=-2.162109375, output=-0.557451608157
			11'd1578: out = 32'b10000000000000000100011111000101; // input=-2.166015625, output=-0.560690352499
			11'd1579: out = 32'b10000000000000000100100000101111; // input=-2.169921875, output=-0.563920541396
			11'd1580: out = 32'b10000000000000000100100010011000; // input=-2.173828125, output=-0.567142125559
			11'd1581: out = 32'b10000000000000000100100100000001; // input=-2.177734375, output=-0.570355055831
			11'd1582: out = 32'b10000000000000000100100101101010; // input=-2.181640625, output=-0.573559283187
			11'd1583: out = 32'b10000000000000000100100111010011; // input=-2.185546875, output=-0.576754758734
			11'd1584: out = 32'b10000000000000000100101000111100; // input=-2.189453125, output=-0.579941433713
			11'd1585: out = 32'b10000000000000000100101010100100; // input=-2.193359375, output=-0.583119259499
			11'd1586: out = 32'b10000000000000000100101100001011; // input=-2.197265625, output=-0.586288187603
			11'd1587: out = 32'b10000000000000000100101101110011; // input=-2.201171875, output=-0.58944816967
			11'd1588: out = 32'b10000000000000000100101111011010; // input=-2.205078125, output=-0.592599157484
			11'd1589: out = 32'b10000000000000000100110001000001; // input=-2.208984375, output=-0.595741102963
			11'd1590: out = 32'b10000000000000000100110010101000; // input=-2.212890625, output=-0.598873958166
			11'd1591: out = 32'b10000000000000000100110100001110; // input=-2.216796875, output=-0.601997675289
			11'd1592: out = 32'b10000000000000000100110101110100; // input=-2.220703125, output=-0.605112206669
			11'd1593: out = 32'b10000000000000000100110111011010; // input=-2.224609375, output=-0.60821750478
			11'd1594: out = 32'b10000000000000000100111001000000; // input=-2.228515625, output=-0.611313522241
			11'd1595: out = 32'b10000000000000000100111010100101; // input=-2.232421875, output=-0.61440021181
			11'd1596: out = 32'b10000000000000000100111100001010; // input=-2.236328125, output=-0.617477526387
			11'd1597: out = 32'b10000000000000000100111101101110; // input=-2.240234375, output=-0.620545419017
			11'd1598: out = 32'b10000000000000000100111111010010; // input=-2.244140625, output=-0.623603842888
			11'd1599: out = 32'b10000000000000000101000000110110; // input=-2.248046875, output=-0.626652751331
			11'd1600: out = 32'b10000000000000000101000010011010; // input=-2.251953125, output=-0.629692097824
			11'd1601: out = 32'b10000000000000000101000011111101; // input=-2.255859375, output=-0.63272183599
			11'd1602: out = 32'b10000000000000000101000101100000; // input=-2.259765625, output=-0.635741919599
			11'd1603: out = 32'b10000000000000000101000111000011; // input=-2.263671875, output=-0.638752302569
			11'd1604: out = 32'b10000000000000000101001000100101; // input=-2.267578125, output=-0.641752938965
			11'd1605: out = 32'b10000000000000000101001010000111; // input=-2.271484375, output=-0.644743783001
			11'd1606: out = 32'b10000000000000000101001011101001; // input=-2.275390625, output=-0.647724789039
			11'd1607: out = 32'b10000000000000000101001101001010; // input=-2.279296875, output=-0.650695911595
			11'd1608: out = 32'b10000000000000000101001110101011; // input=-2.283203125, output=-0.653657105331
			11'd1609: out = 32'b10000000000000000101010000001100; // input=-2.287109375, output=-0.656608325064
			11'd1610: out = 32'b10000000000000000101010001101100; // input=-2.291015625, output=-0.659549525762
			11'd1611: out = 32'b10000000000000000101010011001100; // input=-2.294921875, output=-0.662480662545
			11'd1612: out = 32'b10000000000000000101010100101100; // input=-2.298828125, output=-0.665401690689
			11'd1613: out = 32'b10000000000000000101010110001011; // input=-2.302734375, output=-0.668312565622
			11'd1614: out = 32'b10000000000000000101010111101010; // input=-2.306640625, output=-0.671213242927
			11'd1615: out = 32'b10000000000000000101011001001001; // input=-2.310546875, output=-0.674103678343
			11'd1616: out = 32'b10000000000000000101011010100111; // input=-2.314453125, output=-0.676983827767
			11'd1617: out = 32'b10000000000000000101011100000101; // input=-2.318359375, output=-0.679853647251
			11'd1618: out = 32'b10000000000000000101011101100011; // input=-2.322265625, output=-0.682713093005
			11'd1619: out = 32'b10000000000000000101011111000000; // input=-2.326171875, output=-0.685562121397
			11'd1620: out = 32'b10000000000000000101100000011110; // input=-2.330078125, output=-0.688400688954
			11'd1621: out = 32'b10000000000000000101100001111010; // input=-2.333984375, output=-0.691228752363
			11'd1622: out = 32'b10000000000000000101100011010111; // input=-2.337890625, output=-0.694046268473
			11'd1623: out = 32'b10000000000000000101100100110010; // input=-2.341796875, output=-0.69685319429
			11'd1624: out = 32'b10000000000000000101100110001110; // input=-2.345703125, output=-0.699649486985
			11'd1625: out = 32'b10000000000000000101100111101001; // input=-2.349609375, output=-0.702435103889
			11'd1626: out = 32'b10000000000000000101101001000100; // input=-2.353515625, output=-0.705210002498
			11'd1627: out = 32'b10000000000000000101101010011111; // input=-2.357421875, output=-0.707974140471
			11'd1628: out = 32'b10000000000000000101101011111001; // input=-2.361328125, output=-0.710727475628
			11'd1629: out = 32'b10000000000000000101101101010011; // input=-2.365234375, output=-0.713469965959
			11'd1630: out = 32'b10000000000000000101101110101100; // input=-2.369140625, output=-0.716201569616
			11'd1631: out = 32'b10000000000000000101110000000110; // input=-2.373046875, output=-0.718922244918
			11'd1632: out = 32'b10000000000000000101110001011110; // input=-2.376953125, output=-0.721631950352
			11'd1633: out = 32'b10000000000000000101110010110111; // input=-2.380859375, output=-0.724330644569
			11'd1634: out = 32'b10000000000000000101110100001111; // input=-2.384765625, output=-0.727018286392
			11'd1635: out = 32'b10000000000000000101110101100111; // input=-2.388671875, output=-0.729694834811
			11'd1636: out = 32'b10000000000000000101110110111110; // input=-2.392578125, output=-0.732360248984
			11'd1637: out = 32'b10000000000000000101111000010101; // input=-2.396484375, output=-0.735014488241
			11'd1638: out = 32'b10000000000000000101111001101100; // input=-2.400390625, output=-0.737657512081
			11'd1639: out = 32'b10000000000000000101111011000010; // input=-2.404296875, output=-0.740289280175
			11'd1640: out = 32'b10000000000000000101111100011000; // input=-2.408203125, output=-0.742909752365
			11'd1641: out = 32'b10000000000000000101111101101101; // input=-2.412109375, output=-0.745518888667
			11'd1642: out = 32'b10000000000000000101111111000010; // input=-2.416015625, output=-0.748116649267
			11'd1643: out = 32'b10000000000000000110000000010111; // input=-2.419921875, output=-0.750702994528
			11'd1644: out = 32'b10000000000000000110000001101011; // input=-2.423828125, output=-0.753277884985
			11'd1645: out = 32'b10000000000000000110000010111111; // input=-2.427734375, output=-0.755841281348
			11'd1646: out = 32'b10000000000000000110000100010011; // input=-2.431640625, output=-0.758393144503
			11'd1647: out = 32'b10000000000000000110000101100110; // input=-2.435546875, output=-0.760933435512
			11'd1648: out = 32'b10000000000000000110000110111001; // input=-2.439453125, output=-0.763462115613
			11'd1649: out = 32'b10000000000000000110001000001100; // input=-2.443359375, output=-0.765979146221
			11'd1650: out = 32'b10000000000000000110001001011110; // input=-2.447265625, output=-0.76848448893
			11'd1651: out = 32'b10000000000000000110001010101111; // input=-2.451171875, output=-0.770978105511
			11'd1652: out = 32'b10000000000000000110001100000001; // input=-2.455078125, output=-0.773459957915
			11'd1653: out = 32'b10000000000000000110001101010010; // input=-2.458984375, output=-0.775930008271
			11'd1654: out = 32'b10000000000000000110001110100010; // input=-2.462890625, output=-0.77838821889
			11'd1655: out = 32'b10000000000000000110001111110010; // input=-2.466796875, output=-0.780834552263
			11'd1656: out = 32'b10000000000000000110010001000010; // input=-2.470703125, output=-0.783268971061
			11'd1657: out = 32'b10000000000000000110010010010010; // input=-2.474609375, output=-0.785691438138
			11'd1658: out = 32'b10000000000000000110010011100001; // input=-2.478515625, output=-0.78810191653
			11'd1659: out = 32'b10000000000000000110010100101111; // input=-2.482421875, output=-0.790500369457
			11'd1660: out = 32'b10000000000000000110010101111101; // input=-2.486328125, output=-0.792886760321
			11'd1661: out = 32'b10000000000000000110010111001011; // input=-2.490234375, output=-0.795261052708
			11'd1662: out = 32'b10000000000000000110011000011001; // input=-2.494140625, output=-0.797623210391
			11'd1663: out = 32'b10000000000000000110011001100110; // input=-2.498046875, output=-0.799973197324
			11'd1664: out = 32'b10000000000000000110011010110010; // input=-2.501953125, output=-0.802310977651
			11'd1665: out = 32'b10000000000000000110011011111110; // input=-2.505859375, output=-0.804636515699
			11'd1666: out = 32'b10000000000000000110011101001010; // input=-2.509765625, output=-0.806949775984
			11'd1667: out = 32'b10000000000000000110011110010110; // input=-2.513671875, output=-0.809250723208
			11'd1668: out = 32'b10000000000000000110011111100001; // input=-2.517578125, output=-0.811539322262
			11'd1669: out = 32'b10000000000000000110100000101011; // input=-2.521484375, output=-0.813815538224
			11'd1670: out = 32'b10000000000000000110100001110101; // input=-2.525390625, output=-0.816079336362
			11'd1671: out = 32'b10000000000000000110100010111111; // input=-2.529296875, output=-0.818330682134
			11'd1672: out = 32'b10000000000000000110100100001000; // input=-2.533203125, output=-0.820569541186
			11'd1673: out = 32'b10000000000000000110100101010001; // input=-2.537109375, output=-0.822795879357
			11'd1674: out = 32'b10000000000000000110100110011010; // input=-2.541015625, output=-0.825009662675
			11'd1675: out = 32'b10000000000000000110100111100010; // input=-2.544921875, output=-0.82721085736
			11'd1676: out = 32'b10000000000000000110101000101010; // input=-2.548828125, output=-0.829399429826
			11'd1677: out = 32'b10000000000000000110101001110001; // input=-2.552734375, output=-0.831575346677
			11'd1678: out = 32'b10000000000000000110101010111000; // input=-2.556640625, output=-0.833738574711
			11'd1679: out = 32'b10000000000000000110101011111110; // input=-2.560546875, output=-0.83588908092
			11'd1680: out = 32'b10000000000000000110101101000100; // input=-2.564453125, output=-0.83802683249
			11'd1681: out = 32'b10000000000000000110101110001010; // input=-2.568359375, output=-0.840151796802
			11'd1682: out = 32'b10000000000000000110101111001111; // input=-2.572265625, output=-0.842263941431
			11'd1683: out = 32'b10000000000000000110110000010100; // input=-2.576171875, output=-0.844363234149
			11'd1684: out = 32'b10000000000000000110110001011000; // input=-2.580078125, output=-0.846449642922
			11'd1685: out = 32'b10000000000000000110110010011100; // input=-2.583984375, output=-0.848523135916
			11'd1686: out = 32'b10000000000000000110110011100000; // input=-2.587890625, output=-0.85058368149
			11'd1687: out = 32'b10000000000000000110110100100011; // input=-2.591796875, output=-0.852631248204
			11'd1688: out = 32'b10000000000000000110110101100110; // input=-2.595703125, output=-0.854665804814
			11'd1689: out = 32'b10000000000000000110110110101000; // input=-2.599609375, output=-0.856687320275
			11'd1690: out = 32'b10000000000000000110110111101010; // input=-2.603515625, output=-0.858695763742
			11'd1691: out = 32'b10000000000000000110111000101011; // input=-2.607421875, output=-0.860691104568
			11'd1692: out = 32'b10000000000000000110111001101100; // input=-2.611328125, output=-0.862673312307
			11'd1693: out = 32'b10000000000000000110111010101101; // input=-2.615234375, output=-0.864642356712
			11'd1694: out = 32'b10000000000000000110111011101101; // input=-2.619140625, output=-0.866598207739
			11'd1695: out = 32'b10000000000000000110111100101100; // input=-2.623046875, output=-0.868540835543
			11'd1696: out = 32'b10000000000000000110111101101100; // input=-2.626953125, output=-0.870470210483
			11'd1697: out = 32'b10000000000000000110111110101010; // input=-2.630859375, output=-0.872386303118
			11'd1698: out = 32'b10000000000000000110111111101001; // input=-2.634765625, output=-0.874289084212
			11'd1699: out = 32'b10000000000000000111000000100111; // input=-2.638671875, output=-0.87617852473
			11'd1700: out = 32'b10000000000000000111000001100100; // input=-2.642578125, output=-0.878054595842
			11'd1701: out = 32'b10000000000000000111000010100001; // input=-2.646484375, output=-0.879917268921
			11'd1702: out = 32'b10000000000000000111000011011110; // input=-2.650390625, output=-0.881766515544
			11'd1703: out = 32'b10000000000000000111000100011010; // input=-2.654296875, output=-0.883602307496
			11'd1704: out = 32'b10000000000000000111000101010110; // input=-2.658203125, output=-0.885424616764
			11'd1705: out = 32'b10000000000000000111000110010001; // input=-2.662109375, output=-0.887233415541
			11'd1706: out = 32'b10000000000000000111000111001100; // input=-2.666015625, output=-0.889028676228
			11'd1707: out = 32'b10000000000000000111001000000110; // input=-2.669921875, output=-0.890810371432
			11'd1708: out = 32'b10000000000000000111001001000000; // input=-2.673828125, output=-0.892578473965
			11'd1709: out = 32'b10000000000000000111001001111010; // input=-2.677734375, output=-0.894332956848
			11'd1710: out = 32'b10000000000000000111001010110011; // input=-2.681640625, output=-0.896073793311
			11'd1711: out = 32'b10000000000000000111001011101011; // input=-2.685546875, output=-0.897800956791
			11'd1712: out = 32'b10000000000000000111001100100011; // input=-2.689453125, output=-0.899514420932
			11'd1713: out = 32'b10000000000000000111001101011011; // input=-2.693359375, output=-0.90121415959
			11'd1714: out = 32'b10000000000000000111001110010010; // input=-2.697265625, output=-0.902900146829
			11'd1715: out = 32'b10000000000000000111001111001001; // input=-2.701171875, output=-0.904572356923
			11'd1716: out = 32'b10000000000000000111001111111111; // input=-2.705078125, output=-0.906230764355
			11'd1717: out = 32'b10000000000000000111010000110101; // input=-2.708984375, output=-0.907875343821
			11'd1718: out = 32'b10000000000000000111010001101011; // input=-2.712890625, output=-0.909506070226
			11'd1719: out = 32'b10000000000000000111010010100000; // input=-2.716796875, output=-0.911122918687
			11'd1720: out = 32'b10000000000000000111010011010100; // input=-2.720703125, output=-0.912725864533
			11'd1721: out = 32'b10000000000000000111010100001000; // input=-2.724609375, output=-0.914314883306
			11'd1722: out = 32'b10000000000000000111010100111100; // input=-2.728515625, output=-0.915889950759
			11'd1723: out = 32'b10000000000000000111010101101111; // input=-2.732421875, output=-0.917451042858
			11'd1724: out = 32'b10000000000000000111010110100010; // input=-2.736328125, output=-0.918998135783
			11'd1725: out = 32'b10000000000000000111010111010100; // input=-2.740234375, output=-0.920531205927
			11'd1726: out = 32'b10000000000000000111011000000110; // input=-2.744140625, output=-0.922050229897
			11'd1727: out = 32'b10000000000000000111011000110111; // input=-2.748046875, output=-0.923555184515
			11'd1728: out = 32'b10000000000000000111011001101000; // input=-2.751953125, output=-0.925046046817
			11'd1729: out = 32'b10000000000000000111011010011000; // input=-2.755859375, output=-0.926522794055
			11'd1730: out = 32'b10000000000000000111011011001000; // input=-2.759765625, output=-0.927985403695
			11'd1731: out = 32'b10000000000000000111011011111000; // input=-2.763671875, output=-0.929433853419
			11'd1732: out = 32'b10000000000000000111011100100111; // input=-2.767578125, output=-0.930868121127
			11'd1733: out = 32'b10000000000000000111011101010101; // input=-2.771484375, output=-0.932288184932
			11'd1734: out = 32'b10000000000000000111011110000011; // input=-2.775390625, output=-0.933694023166
			11'd1735: out = 32'b10000000000000000111011110110001; // input=-2.779296875, output=-0.935085614378
			11'd1736: out = 32'b10000000000000000111011111011110; // input=-2.783203125, output=-0.936462937335
			11'd1737: out = 32'b10000000000000000111100000001011; // input=-2.787109375, output=-0.937825971019
			11'd1738: out = 32'b10000000000000000111100000110111; // input=-2.791015625, output=-0.939174694632
			11'd1739: out = 32'b10000000000000000111100001100011; // input=-2.794921875, output=-0.940509087596
			11'd1740: out = 32'b10000000000000000111100010001110; // input=-2.798828125, output=-0.941829129547
			11'd1741: out = 32'b10000000000000000111100010111001; // input=-2.802734375, output=-0.943134800345
			11'd1742: out = 32'b10000000000000000111100011100011; // input=-2.806640625, output=-0.944426080067
			11'd1743: out = 32'b10000000000000000111100100001101; // input=-2.810546875, output=-0.945702949008
			11'd1744: out = 32'b10000000000000000111100100110110; // input=-2.814453125, output=-0.946965387686
			11'd1745: out = 32'b10000000000000000111100101011111; // input=-2.818359375, output=-0.948213376837
			11'd1746: out = 32'b10000000000000000111100110000111; // input=-2.822265625, output=-0.949446897419
			11'd1747: out = 32'b10000000000000000111100110101111; // input=-2.826171875, output=-0.950665930609
			11'd1748: out = 32'b10000000000000000111100111010111; // input=-2.830078125, output=-0.951870457806
			11'd1749: out = 32'b10000000000000000111100111111110; // input=-2.833984375, output=-0.953060460632
			11'd1750: out = 32'b10000000000000000111101000100100; // input=-2.837890625, output=-0.954235920927
			11'd1751: out = 32'b10000000000000000111101001001010; // input=-2.841796875, output=-0.955396820757
			11'd1752: out = 32'b10000000000000000111101001110000; // input=-2.845703125, output=-0.956543142406
			11'd1753: out = 32'b10000000000000000111101010010101; // input=-2.849609375, output=-0.957674868384
			11'd1754: out = 32'b10000000000000000111101010111010; // input=-2.853515625, output=-0.958791981422
			11'd1755: out = 32'b10000000000000000111101011011110; // input=-2.857421875, output=-0.959894464473
			11'd1756: out = 32'b10000000000000000111101100000001; // input=-2.861328125, output=-0.960982300717
			11'd1757: out = 32'b10000000000000000111101100100101; // input=-2.865234375, output=-0.962055473552
			11'd1758: out = 32'b10000000000000000111101101000111; // input=-2.869140625, output=-0.963113966605
			11'd1759: out = 32'b10000000000000000111101101101010; // input=-2.873046875, output=-0.964157763723
			11'd1760: out = 32'b10000000000000000111101110001011; // input=-2.876953125, output=-0.965186848981
			11'd1761: out = 32'b10000000000000000111101110101100; // input=-2.880859375, output=-0.966201206674
			11'd1762: out = 32'b10000000000000000111101111001101; // input=-2.884765625, output=-0.967200821326
			11'd1763: out = 32'b10000000000000000111101111101110; // input=-2.888671875, output=-0.968185677683
			11'd1764: out = 32'b10000000000000000111110000001101; // input=-2.892578125, output=-0.969155760718
			11'd1765: out = 32'b10000000000000000111110000101101; // input=-2.896484375, output=-0.970111055629
			11'd1766: out = 32'b10000000000000000111110001001011; // input=-2.900390625, output=-0.971051547838
			11'd1767: out = 32'b10000000000000000111110001101010; // input=-2.904296875, output=-0.971977222996
			11'd1768: out = 32'b10000000000000000111110010001000; // input=-2.908203125, output=-0.972888066977
			11'd1769: out = 32'b10000000000000000111110010100101; // input=-2.912109375, output=-0.973784065883
			11'd1770: out = 32'b10000000000000000111110011000010; // input=-2.916015625, output=-0.974665206042
			11'd1771: out = 32'b10000000000000000111110011011110; // input=-2.919921875, output=-0.975531474009
			11'd1772: out = 32'b10000000000000000111110011111010; // input=-2.923828125, output=-0.976382856567
			11'd1773: out = 32'b10000000000000000111110100010110; // input=-2.927734375, output=-0.977219340723
			11'd1774: out = 32'b10000000000000000111110100110000; // input=-2.931640625, output=-0.978040913714
			11'd1775: out = 32'b10000000000000000111110101001011; // input=-2.935546875, output=-0.978847563005
			11'd1776: out = 32'b10000000000000000111110101100101; // input=-2.939453125, output=-0.979639276285
			11'd1777: out = 32'b10000000000000000111110101111110; // input=-2.943359375, output=-0.980416041476
			11'd1778: out = 32'b10000000000000000111110110010111; // input=-2.947265625, output=-0.981177846724
			11'd1779: out = 32'b10000000000000000111110110110000; // input=-2.951171875, output=-0.981924680406
			11'd1780: out = 32'b10000000000000000111110111001000; // input=-2.955078125, output=-0.982656531125
			11'd1781: out = 32'b10000000000000000111110111011111; // input=-2.958984375, output=-0.983373387714
			11'd1782: out = 32'b10000000000000000111110111110110; // input=-2.962890625, output=-0.984075239235
			11'd1783: out = 32'b10000000000000000111111000001101; // input=-2.966796875, output=-0.984762074979
			11'd1784: out = 32'b10000000000000000111111000100011; // input=-2.970703125, output=-0.985433884466
			11'd1785: out = 32'b10000000000000000111111000111000; // input=-2.974609375, output=-0.986090657443
			11'd1786: out = 32'b10000000000000000111111001001101; // input=-2.978515625, output=-0.986732383891
			11'd1787: out = 32'b10000000000000000111111001100010; // input=-2.982421875, output=-0.987359054016
			11'd1788: out = 32'b10000000000000000111111001110110; // input=-2.986328125, output=-0.987970658257
			11'd1789: out = 32'b10000000000000000111111010001001; // input=-2.990234375, output=-0.988567187281
			11'd1790: out = 32'b10000000000000000111111010011100; // input=-2.994140625, output=-0.989148631986
			11'd1791: out = 32'b10000000000000000111111010101111; // input=-2.998046875, output=-0.9897149835
			11'd1792: out = 32'b10000000000000000111111011000001; // input=-3.001953125, output=-0.990266233181
			11'd1793: out = 32'b10000000000000000111111011010011; // input=-3.005859375, output=-0.990802372617
			11'd1794: out = 32'b10000000000000000111111011100100; // input=-3.009765625, output=-0.991323393629
			11'd1795: out = 32'b10000000000000000111111011110100; // input=-3.013671875, output=-0.991829288265
			11'd1796: out = 32'b10000000000000000111111100000100; // input=-3.017578125, output=-0.992320048806
			11'd1797: out = 32'b10000000000000000111111100010100; // input=-3.021484375, output=-0.992795667765
			11'd1798: out = 32'b10000000000000000111111100100011; // input=-3.025390625, output=-0.993256137883
			11'd1799: out = 32'b10000000000000000111111100110010; // input=-3.029296875, output=-0.993701452134
			11'd1800: out = 32'b10000000000000000111111101000000; // input=-3.033203125, output=-0.994131603724
			11'd1801: out = 32'b10000000000000000111111101001101; // input=-3.037109375, output=-0.994546586089
			11'd1802: out = 32'b10000000000000000111111101011010; // input=-3.041015625, output=-0.994946392896
			11'd1803: out = 32'b10000000000000000111111101100111; // input=-3.044921875, output=-0.995331018046
			11'd1804: out = 32'b10000000000000000111111101110011; // input=-3.048828125, output=-0.995700455669
			11'd1805: out = 32'b10000000000000000111111101111111; // input=-3.052734375, output=-0.996054700128
			11'd1806: out = 32'b10000000000000000111111110001010; // input=-3.056640625, output=-0.996393746017
			11'd1807: out = 32'b10000000000000000111111110010100; // input=-3.060546875, output=-0.996717588164
			11'd1808: out = 32'b10000000000000000111111110011111; // input=-3.064453125, output=-0.997026221627
			11'd1809: out = 32'b10000000000000000111111110101000; // input=-3.068359375, output=-0.997319641697
			11'd1810: out = 32'b10000000000000000111111110110001; // input=-3.072265625, output=-0.997597843896
			11'd1811: out = 32'b10000000000000000111111110111010; // input=-3.076171875, output=-0.997860823979
			11'd1812: out = 32'b10000000000000000111111111000010; // input=-3.080078125, output=-0.998108577933
			11'd1813: out = 32'b10000000000000000111111111001010; // input=-3.083984375, output=-0.998341101979
			11'd1814: out = 32'b10000000000000000111111111010001; // input=-3.087890625, output=-0.998558392568
			11'd1815: out = 32'b10000000000000000111111111010111; // input=-3.091796875, output=-0.998760446384
			11'd1816: out = 32'b10000000000000000111111111011110; // input=-3.095703125, output=-0.998947260345
			11'd1817: out = 32'b10000000000000000111111111100011; // input=-3.099609375, output=-0.999118831599
			11'd1818: out = 32'b10000000000000000111111111101000; // input=-3.103515625, output=-0.99927515753
			11'd1819: out = 32'b10000000000000000111111111101101; // input=-3.107421875, output=-0.999416235751
			11'd1820: out = 32'b10000000000000000111111111110001; // input=-3.111328125, output=-0.99954206411
			11'd1821: out = 32'b10000000000000000111111111110101; // input=-3.115234375, output=-0.999652640687
			11'd1822: out = 32'b10000000000000000111111111111000; // input=-3.119140625, output=-0.999747963794
			11'd1823: out = 32'b10000000000000000111111111111010; // input=-3.123046875, output=-0.999828031977
			11'd1824: out = 32'b10000000000000000111111111111100; // input=-3.126953125, output=-0.999892844015
			11'd1825: out = 32'b10000000000000000111111111111110; // input=-3.130859375, output=-0.999942398918
			11'd1826: out = 32'b10000000000000000111111111111111; // input=-3.134765625, output=-0.999976695931
			11'd1827: out = 32'b10000000000000000111111111111111; // input=-3.138671875, output=-0.999995734529
			11'd1828: out = 32'b10000000000000000111111111111111; // input=-3.142578125, output=-0.999999514423
			11'd1829: out = 32'b10000000000000000111111111111111; // input=-3.146484375, output=-0.999988035555
			11'd1830: out = 32'b10000000000000000111111111111111; // input=-3.150390625, output=-0.999961298099
			11'd1831: out = 32'b10000000000000000111111111111101; // input=-3.154296875, output=-0.999919302465
			11'd1832: out = 32'b10000000000000000111111111111011; // input=-3.158203125, output=-0.999862049292
			11'd1833: out = 32'b10000000000000000111111111111001; // input=-3.162109375, output=-0.999789539454
			11'd1834: out = 32'b10000000000000000111111111110110; // input=-3.166015625, output=-0.999701774058
			11'd1835: out = 32'b10000000000000000111111111110011; // input=-3.169921875, output=-0.999598754443
			11'd1836: out = 32'b10000000000000000111111111101111; // input=-3.173828125, output=-0.999480482181
			11'd1837: out = 32'b10000000000000000111111111101011; // input=-3.177734375, output=-0.999346959076
			11'd1838: out = 32'b10000000000000000111111111100110; // input=-3.181640625, output=-0.999198187167
			11'd1839: out = 32'b10000000000000000111111111100000; // input=-3.185546875, output=-0.999034168722
			11'd1840: out = 32'b10000000000000000111111111011010; // input=-3.189453125, output=-0.998854906245
			11'd1841: out = 32'b10000000000000000111111111010100; // input=-3.193359375, output=-0.998660402471
			11'd1842: out = 32'b10000000000000000111111111001101; // input=-3.197265625, output=-0.998450660368
			11'd1843: out = 32'b10000000000000000111111111000110; // input=-3.201171875, output=-0.998225683137
			11'd1844: out = 32'b10000000000000000111111110111110; // input=-3.205078125, output=-0.997985474209
			11'd1845: out = 32'b10000000000000000111111110110110; // input=-3.208984375, output=-0.997730037251
			11'd1846: out = 32'b10000000000000000111111110101101; // input=-3.212890625, output=-0.997459376161
			11'd1847: out = 32'b10000000000000000111111110100011; // input=-3.216796875, output=-0.997173495067
			11'd1848: out = 32'b10000000000000000111111110011010; // input=-3.220703125, output=-0.996872398333
			11'd1849: out = 32'b10000000000000000111111110001111; // input=-3.224609375, output=-0.996556090553
			11'd1850: out = 32'b10000000000000000111111110000100; // input=-3.228515625, output=-0.996224576552
			11'd1851: out = 32'b10000000000000000111111101111001; // input=-3.232421875, output=-0.995877861391
			11'd1852: out = 32'b10000000000000000111111101101101; // input=-3.236328125, output=-0.995515950358
			11'd1853: out = 32'b10000000000000000111111101100001; // input=-3.240234375, output=-0.995138848977
			11'd1854: out = 32'b10000000000000000111111101010100; // input=-3.244140625, output=-0.994746563001
			11'd1855: out = 32'b10000000000000000111111101000111; // input=-3.248046875, output=-0.994339098417
			11'd1856: out = 32'b10000000000000000111111100111001; // input=-3.251953125, output=-0.993916461441
			11'd1857: out = 32'b10000000000000000111111100101010; // input=-3.255859375, output=-0.993478658524
			11'd1858: out = 32'b10000000000000000111111100011011; // input=-3.259765625, output=-0.993025696344
			11'd1859: out = 32'b10000000000000000111111100001100; // input=-3.263671875, output=-0.992557581813
			11'd1860: out = 32'b10000000000000000111111011111100; // input=-3.267578125, output=-0.992074322076
			11'd1861: out = 32'b10000000000000000111111011101100; // input=-3.271484375, output=-0.991575924504
			11'd1862: out = 32'b10000000000000000111111011011011; // input=-3.275390625, output=-0.991062396704
			11'd1863: out = 32'b10000000000000000111111011001010; // input=-3.279296875, output=-0.990533746511
			11'd1864: out = 32'b10000000000000000111111010111000; // input=-3.283203125, output=-0.989989981992
			11'd1865: out = 32'b10000000000000000111111010100110; // input=-3.287109375, output=-0.989431111444
			11'd1866: out = 32'b10000000000000000111111010010011; // input=-3.291015625, output=-0.988857143395
			11'd1867: out = 32'b10000000000000000111111010000000; // input=-3.294921875, output=-0.988268086602
			11'd1868: out = 32'b10000000000000000111111001101100; // input=-3.298828125, output=-0.987663950053
			11'd1869: out = 32'b10000000000000000111111001010111; // input=-3.302734375, output=-0.987044742969
			11'd1870: out = 32'b10000000000000000111111001000011; // input=-3.306640625, output=-0.986410474795
			11'd1871: out = 32'b10000000000000000111111000101101; // input=-3.310546875, output=-0.985761155212
			11'd1872: out = 32'b10000000000000000111111000011000; // input=-3.314453125, output=-0.985096794126
			11'd1873: out = 32'b10000000000000000111111000000001; // input=-3.318359375, output=-0.984417401675
			11'd1874: out = 32'b10000000000000000111110111101011; // input=-3.322265625, output=-0.983722988226
			11'd1875: out = 32'b10000000000000000111110111010011; // input=-3.326171875, output=-0.983013564374
			11'd1876: out = 32'b10000000000000000111110110111100; // input=-3.330078125, output=-0.982289140945
			11'd1877: out = 32'b10000000000000000111110110100011; // input=-3.333984375, output=-0.981549728992
			11'd1878: out = 32'b10000000000000000111110110001011; // input=-3.337890625, output=-0.980795339798
			11'd1879: out = 32'b10000000000000000111110101110001; // input=-3.341796875, output=-0.980025984873
			11'd1880: out = 32'b10000000000000000111110101011000; // input=-3.345703125, output=-0.979241675958
			11'd1881: out = 32'b10000000000000000111110100111110; // input=-3.349609375, output=-0.978442425019
			11'd1882: out = 32'b10000000000000000111110100100011; // input=-3.353515625, output=-0.977628244254
			11'd1883: out = 32'b10000000000000000111110100001000; // input=-3.357421875, output=-0.976799146083
			11'd1884: out = 32'b10000000000000000111110011101100; // input=-3.361328125, output=-0.97595514316
			11'd1885: out = 32'b10000000000000000111110011010000; // input=-3.365234375, output=-0.975096248362
			11'd1886: out = 32'b10000000000000000111110010110011; // input=-3.369140625, output=-0.974222474795
			11'd1887: out = 32'b10000000000000000111110010010110; // input=-3.373046875, output=-0.973333835791
			11'd1888: out = 32'b10000000000000000111110001111001; // input=-3.376953125, output=-0.972430344911
			11'd1889: out = 32'b10000000000000000111110001011011; // input=-3.380859375, output=-0.97151201594
			11'd1890: out = 32'b10000000000000000111110000111100; // input=-3.384765625, output=-0.970578862891
			11'd1891: out = 32'b10000000000000000111110000011101; // input=-3.388671875, output=-0.969630900003
			11'd1892: out = 32'b10000000000000000111101111111101; // input=-3.392578125, output=-0.96866814174
			11'd1893: out = 32'b10000000000000000111101111011101; // input=-3.396484375, output=-0.967690602793
			11'd1894: out = 32'b10000000000000000111101110111101; // input=-3.400390625, output=-0.966698298078
			11'd1895: out = 32'b10000000000000000111101110011100; // input=-3.404296875, output=-0.965691242737
			11'd1896: out = 32'b10000000000000000111101101111010; // input=-3.408203125, output=-0.964669452135
			11'd1897: out = 32'b10000000000000000111101101011000; // input=-3.412109375, output=-0.963632941864
			11'd1898: out = 32'b10000000000000000111101100110110; // input=-3.416015625, output=-0.96258172774
			11'd1899: out = 32'b10000000000000000111101100010011; // input=-3.419921875, output=-0.961515825803
			11'd1900: out = 32'b10000000000000000111101011110000; // input=-3.423828125, output=-0.960435252318
			11'd1901: out = 32'b10000000000000000111101011001100; // input=-3.427734375, output=-0.959340023773
			11'd1902: out = 32'b10000000000000000111101010100111; // input=-3.431640625, output=-0.958230156879
			11'd1903: out = 32'b10000000000000000111101010000010; // input=-3.435546875, output=-0.957105668571
			11'd1904: out = 32'b10000000000000000111101001011101; // input=-3.439453125, output=-0.955966576009
			11'd1905: out = 32'b10000000000000000111101000110111; // input=-3.443359375, output=-0.954812896573
			11'd1906: out = 32'b10000000000000000111101000010001; // input=-3.447265625, output=-0.953644647867
			11'd1907: out = 32'b10000000000000000111100111101010; // input=-3.451171875, output=-0.952461847717
			11'd1908: out = 32'b10000000000000000111100111000011; // input=-3.455078125, output=-0.951264514171
			11'd1909: out = 32'b10000000000000000111100110011011; // input=-3.458984375, output=-0.950052665499
			11'd1910: out = 32'b10000000000000000111100101110011; // input=-3.462890625, output=-0.948826320192
			11'd1911: out = 32'b10000000000000000111100101001010; // input=-3.466796875, output=-0.947585496963
			11'd1912: out = 32'b10000000000000000111100100100001; // input=-3.470703125, output=-0.946330214745
			11'd1913: out = 32'b10000000000000000111100011111000; // input=-3.474609375, output=-0.945060492692
			11'd1914: out = 32'b10000000000000000111100011001110; // input=-3.478515625, output=-0.943776350179
			11'd1915: out = 32'b10000000000000000111100010100011; // input=-3.482421875, output=-0.9424778068
			11'd1916: out = 32'b10000000000000000111100001111000; // input=-3.486328125, output=-0.94116488237
			11'd1917: out = 32'b10000000000000000111100001001101; // input=-3.490234375, output=-0.939837596921
			11'd1918: out = 32'b10000000000000000111100000100001; // input=-3.494140625, output=-0.938495970706
			11'd1919: out = 32'b10000000000000000111011111110100; // input=-3.498046875, output=-0.937140024198
			11'd1920: out = 32'b10000000000000000111011111000111; // input=-3.501953125, output=-0.935769778086
			11'd1921: out = 32'b10000000000000000111011110011010; // input=-3.505859375, output=-0.934385253279
			11'd1922: out = 32'b10000000000000000111011101101100; // input=-3.509765625, output=-0.932986470902
			11'd1923: out = 32'b10000000000000000111011100111110; // input=-3.513671875, output=-0.931573452299
			11'd1924: out = 32'b10000000000000000111011100001111; // input=-3.517578125, output=-0.930146219032
			11'd1925: out = 32'b10000000000000000111011011100000; // input=-3.521484375, output=-0.928704792878
			11'd1926: out = 32'b10000000000000000111011010110000; // input=-3.525390625, output=-0.927249195831
			11'd1927: out = 32'b10000000000000000111011010000000; // input=-3.529296875, output=-0.925779450103
			11'd1928: out = 32'b10000000000000000111011001001111; // input=-3.533203125, output=-0.924295578119
			11'd1929: out = 32'b10000000000000000111011000011110; // input=-3.537109375, output=-0.922797602521
			11'd1930: out = 32'b10000000000000000111010111101101; // input=-3.541015625, output=-0.921285546168
			11'd1931: out = 32'b10000000000000000111010110111011; // input=-3.544921875, output=-0.919759432131
			11'd1932: out = 32'b10000000000000000111010110001000; // input=-3.548828125, output=-0.918219283696
			11'd1933: out = 32'b10000000000000000111010101010101; // input=-3.552734375, output=-0.916665124365
			11'd1934: out = 32'b10000000000000000111010100100010; // input=-3.556640625, output=-0.915096977852
			11'd1935: out = 32'b10000000000000000111010011101110; // input=-3.560546875, output=-0.913514868085
			11'd1936: out = 32'b10000000000000000111010010111010; // input=-3.564453125, output=-0.911918819205
			11'd1937: out = 32'b10000000000000000111010010000101; // input=-3.568359375, output=-0.910308855566
			11'd1938: out = 32'b10000000000000000111010001010000; // input=-3.572265625, output=-0.908685001733
			11'd1939: out = 32'b10000000000000000111010000011010; // input=-3.576171875, output=-0.907047282486
			11'd1940: out = 32'b10000000000000000111001111100100; // input=-3.580078125, output=-0.905395722813
			11'd1941: out = 32'b10000000000000000111001110101101; // input=-3.583984375, output=-0.903730347915
			11'd1942: out = 32'b10000000000000000111001101110110; // input=-3.587890625, output=-0.902051183204
			11'd1943: out = 32'b10000000000000000111001100111111; // input=-3.591796875, output=-0.900358254301
			11'd1944: out = 32'b10000000000000000111001100000111; // input=-3.595703125, output=-0.89865158704
			11'd1945: out = 32'b10000000000000000111001011001111; // input=-3.599609375, output=-0.896931207461
			11'd1946: out = 32'b10000000000000000111001010010110; // input=-3.603515625, output=-0.895197141815
			11'd1947: out = 32'b10000000000000000111001001011101; // input=-3.607421875, output=-0.893449416562
			11'd1948: out = 32'b10000000000000000111001000100011; // input=-3.611328125, output=-0.89168805837
			11'd1949: out = 32'b10000000000000000111000111101001; // input=-3.615234375, output=-0.889913094116
			11'd1950: out = 32'b10000000000000000111000110101110; // input=-3.619140625, output=-0.888124550883
			11'd1951: out = 32'b10000000000000000111000101110011; // input=-3.623046875, output=-0.886322455962
			11'd1952: out = 32'b10000000000000000111000100111000; // input=-3.626953125, output=-0.88450683685
			11'd1953: out = 32'b10000000000000000111000011111100; // input=-3.630859375, output=-0.882677721253
			11'd1954: out = 32'b10000000000000000111000010111111; // input=-3.634765625, output=-0.880835137079
			11'd1955: out = 32'b10000000000000000111000010000010; // input=-3.638671875, output=-0.878979112445
			11'd1956: out = 32'b10000000000000000111000001000101; // input=-3.642578125, output=-0.877109675671
			11'd1957: out = 32'b10000000000000000111000000000111; // input=-3.646484375, output=-0.875226855283
			11'd1958: out = 32'b10000000000000000110111111001001; // input=-3.650390625, output=-0.87333068001
			11'd1959: out = 32'b10000000000000000110111110001011; // input=-3.654296875, output=-0.871421178785
			11'd1960: out = 32'b10000000000000000110111101001100; // input=-3.658203125, output=-0.869498380745
			11'd1961: out = 32'b10000000000000000110111100001100; // input=-3.662109375, output=-0.867562315229
			11'd1962: out = 32'b10000000000000000110111011001100; // input=-3.666015625, output=-0.86561301178
			11'd1963: out = 32'b10000000000000000110111010001100; // input=-3.669921875, output=-0.863650500142
			11'd1964: out = 32'b10000000000000000110111001001011; // input=-3.673828125, output=-0.861674810259
			11'd1965: out = 32'b10000000000000000110111000001010; // input=-3.677734375, output=-0.859685972279
			11'd1966: out = 32'b10000000000000000110110111001001; // input=-3.681640625, output=-0.857684016548
			11'd1967: out = 32'b10000000000000000110110110000111; // input=-3.685546875, output=-0.855668973615
			11'd1968: out = 32'b10000000000000000110110101000100; // input=-3.689453125, output=-0.853640874226
			11'd1969: out = 32'b10000000000000000110110100000001; // input=-3.693359375, output=-0.851599749328
			11'd1970: out = 32'b10000000000000000110110010111110; // input=-3.697265625, output=-0.849545630065
			11'd1971: out = 32'b10000000000000000110110001111010; // input=-3.701171875, output=-0.847478547781
			11'd1972: out = 32'b10000000000000000110110000110110; // input=-3.705078125, output=-0.845398534017
			11'd1973: out = 32'b10000000000000000110101111110001; // input=-3.708984375, output=-0.843305620512
			11'd1974: out = 32'b10000000000000000110101110101100; // input=-3.712890625, output=-0.8411998392
			11'd1975: out = 32'b10000000000000000110101101100111; // input=-3.716796875, output=-0.839081222214
			11'd1976: out = 32'b10000000000000000110101100100001; // input=-3.720703125, output=-0.83694980188
			11'd1977: out = 32'b10000000000000000110101011011011; // input=-3.724609375, output=-0.834805610723
			11'd1978: out = 32'b10000000000000000110101010010100; // input=-3.728515625, output=-0.832648681459
			11'd1979: out = 32'b10000000000000000110101001001101; // input=-3.732421875, output=-0.830479047
			11'd1980: out = 32'b10000000000000000110101000000110; // input=-3.736328125, output=-0.828296740453
			11'd1981: out = 32'b10000000000000000110100110111110; // input=-3.740234375, output=-0.826101795117
			11'd1982: out = 32'b10000000000000000110100101110101; // input=-3.744140625, output=-0.823894244484
			11'd1983: out = 32'b10000000000000000110100100101101; // input=-3.748046875, output=-0.821674122238
			11'd1984: out = 32'b10000000000000000110100011100011; // input=-3.751953125, output=-0.819441462256
			11'd1985: out = 32'b10000000000000000110100010011010; // input=-3.755859375, output=-0.817196298606
			11'd1986: out = 32'b10000000000000000110100001010000; // input=-3.759765625, output=-0.814938665546
			11'd1987: out = 32'b10000000000000000110100000000110; // input=-3.763671875, output=-0.812668597524
			11'd1988: out = 32'b10000000000000000110011110111011; // input=-3.767578125, output=-0.810386129179
			11'd1989: out = 32'b10000000000000000110011101110000; // input=-3.771484375, output=-0.808091295339
			11'd1990: out = 32'b10000000000000000110011100100100; // input=-3.775390625, output=-0.80578413102
			11'd1991: out = 32'b10000000000000000110011011011000; // input=-3.779296875, output=-0.803464671426
			11'd1992: out = 32'b10000000000000000110011010001100; // input=-3.783203125, output=-0.801132951951
			11'd1993: out = 32'b10000000000000000110011000111111; // input=-3.787109375, output=-0.798789008172
			11'd1994: out = 32'b10000000000000000110010111110010; // input=-3.791015625, output=-0.796432875855
			11'd1995: out = 32'b10000000000000000110010110100100; // input=-3.794921875, output=-0.794064590953
			11'd1996: out = 32'b10000000000000000110010101010110; // input=-3.798828125, output=-0.791684189602
			11'd1997: out = 32'b10000000000000000110010100001000; // input=-3.802734375, output=-0.789291708124
			11'd1998: out = 32'b10000000000000000110010010111001; // input=-3.806640625, output=-0.786887183026
			11'd1999: out = 32'b10000000000000000110010001101010; // input=-3.810546875, output=-0.784470650998
			11'd2000: out = 32'b10000000000000000110010000011010; // input=-3.814453125, output=-0.782042148913
			11'd2001: out = 32'b10000000000000000110001111001010; // input=-3.818359375, output=-0.779601713826
			11'd2002: out = 32'b10000000000000000110001101111010; // input=-3.822265625, output=-0.777149382977
			11'd2003: out = 32'b10000000000000000110001100101001; // input=-3.826171875, output=-0.774685193784
			11'd2004: out = 32'b10000000000000000110001011011000; // input=-3.830078125, output=-0.772209183849
			11'd2005: out = 32'b10000000000000000110001010000110; // input=-3.833984375, output=-0.769721390951
			11'd2006: out = 32'b10000000000000000110001000110100; // input=-3.837890625, output=-0.767221853052
			11'd2007: out = 32'b10000000000000000110000111100010; // input=-3.841796875, output=-0.764710608291
			11'd2008: out = 32'b10000000000000000110000110001111; // input=-3.845703125, output=-0.762187694988
			11'd2009: out = 32'b10000000000000000110000100111100; // input=-3.849609375, output=-0.759653151638
			11'd2010: out = 32'b10000000000000000110000011101001; // input=-3.853515625, output=-0.757107016915
			11'd2011: out = 32'b10000000000000000110000010010101; // input=-3.857421875, output=-0.754549329671
			11'd2012: out = 32'b10000000000000000110000001000001; // input=-3.861328125, output=-0.751980128932
			11'd2013: out = 32'b10000000000000000101111111101100; // input=-3.865234375, output=-0.749399453902
			11'd2014: out = 32'b10000000000000000101111110010111; // input=-3.869140625, output=-0.746807343958
			11'd2015: out = 32'b10000000000000000101111101000010; // input=-3.873046875, output=-0.744203838653
			11'd2016: out = 32'b10000000000000000101111011101100; // input=-3.876953125, output=-0.741588977713
			11'd2017: out = 32'b10000000000000000101111010010110; // input=-3.880859375, output=-0.738962801038
			11'd2018: out = 32'b10000000000000000101111001000000; // input=-3.884765625, output=-0.736325348699
			11'd2019: out = 32'b10000000000000000101110111101001; // input=-3.888671875, output=-0.733676660942
			11'd2020: out = 32'b10000000000000000101110110010010; // input=-3.892578125, output=-0.731016778181
			11'd2021: out = 32'b10000000000000000101110100111010; // input=-3.896484375, output=-0.728345741004
			11'd2022: out = 32'b10000000000000000101110011100011; // input=-3.900390625, output=-0.725663590167
			11'd2023: out = 32'b10000000000000000101110010001010; // input=-3.904296875, output=-0.722970366596
			11'd2024: out = 32'b10000000000000000101110000110010; // input=-3.908203125, output=-0.720266111387
			11'd2025: out = 32'b10000000000000000101101111011001; // input=-3.912109375, output=-0.717550865803
			11'd2026: out = 32'b10000000000000000101101101111111; // input=-3.916015625, output=-0.714824671276
			11'd2027: out = 32'b10000000000000000101101100100110; // input=-3.919921875, output=-0.712087569404
			11'd2028: out = 32'b10000000000000000101101011001100; // input=-3.923828125, output=-0.709339601952
			11'd2029: out = 32'b10000000000000000101101001110001; // input=-3.927734375, output=-0.70658081085
			11'd2030: out = 32'b10000000000000000101101000010110; // input=-3.931640625, output=-0.703811238194
			11'd2031: out = 32'b10000000000000000101100110111011; // input=-3.935546875, output=-0.701030926245
			11'd2032: out = 32'b10000000000000000101100101100000; // input=-3.939453125, output=-0.698239917426
			11'd2033: out = 32'b10000000000000000101100100000100; // input=-3.943359375, output=-0.695438254325
			11'd2034: out = 32'b10000000000000000101100010101000; // input=-3.947265625, output=-0.692625979692
			11'd2035: out = 32'b10000000000000000101100001001011; // input=-3.951171875, output=-0.689803136439
			11'd2036: out = 32'b10000000000000000101011111101111; // input=-3.955078125, output=-0.686969767639
			11'd2037: out = 32'b10000000000000000101011110010001; // input=-3.958984375, output=-0.684125916525
			11'd2038: out = 32'b10000000000000000101011100110100; // input=-3.962890625, output=-0.681271626491
			11'd2039: out = 32'b10000000000000000101011011010110; // input=-3.966796875, output=-0.678406941091
			11'd2040: out = 32'b10000000000000000101011001111000; // input=-3.970703125, output=-0.675531904035
			11'd2041: out = 32'b10000000000000000101011000011001; // input=-3.974609375, output=-0.672646559194
			11'd2042: out = 32'b10000000000000000101010110111010; // input=-3.978515625, output=-0.669750950593
			11'd2043: out = 32'b10000000000000000101010101011011; // input=-3.982421875, output=-0.666845122418
			11'd2044: out = 32'b10000000000000000101010011111100; // input=-3.986328125, output=-0.663929119006
			11'd2045: out = 32'b10000000000000000101010010011100; // input=-3.990234375, output=-0.661002984852
			11'd2046: out = 32'b10000000000000000101010000111100; // input=-3.994140625, output=-0.658066764607
			11'd2047: out = 32'b10000000000000000101001111011011; // input=-3.998046875, output=-0.655120503072
		endcase
	end
	converter U0 (a, index);

endmodule

module sin_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000000000000001000000; // input=0.001953125, output=0.00195312375824
			11'd1: out = 32'b00000000000000000000000011000000; // input=0.005859375, output=0.00585934147244
			11'd2: out = 32'b00000000000000000000000101000000; // input=0.009765625, output=0.00976546978031
			11'd3: out = 32'b00000000000000000000000111000000; // input=0.013671875, output=0.0136714490791
			11'd4: out = 32'b00000000000000000000001001000000; // input=0.017578125, output=0.0175772197684
			11'd5: out = 32'b00000000000000000000001011000000; // input=0.021484375, output=0.021482722251
			11'd6: out = 32'b00000000000000000000001101000000; // input=0.025390625, output=0.0253878969337
			11'd7: out = 32'b00000000000000000000001111000000; // input=0.029296875, output=0.0292926842283
			11'd8: out = 32'b00000000000000000000010001000000; // input=0.033203125, output=0.0331970245525
			11'd9: out = 32'b00000000000000000000010011000000; // input=0.037109375, output=0.0371008583311
			11'd10: out = 32'b00000000000000000000010101000000; // input=0.041015625, output=0.0410041259961
			11'd11: out = 32'b00000000000000000000010111000000; // input=0.044921875, output=0.0449067679887
			11'd12: out = 32'b00000000000000000000011000111111; // input=0.048828125, output=0.0488087247592
			11'd13: out = 32'b00000000000000000000011010111111; // input=0.052734375, output=0.0527099367686
			11'd14: out = 32'b00000000000000000000011100111111; // input=0.056640625, output=0.0566103444893
			11'd15: out = 32'b00000000000000000000011110111111; // input=0.060546875, output=0.0605098884057
			11'd16: out = 32'b00000000000000000000100000111111; // input=0.064453125, output=0.0644085090157
			11'd17: out = 32'b00000000000000000000100010111110; // input=0.068359375, output=0.0683061468311
			11'd18: out = 32'b00000000000000000000100100111110; // input=0.072265625, output=0.0722027423787
			11'd19: out = 32'b00000000000000000000100110111110; // input=0.076171875, output=0.0760982362014
			11'd20: out = 32'b00000000000000000000101000111101; // input=0.080078125, output=0.0799925688585
			11'd21: out = 32'b00000000000000000000101010111101; // input=0.083984375, output=0.0838856809275
			11'd22: out = 32'b00000000000000000000101100111100; // input=0.087890625, output=0.0877775130042
			11'd23: out = 32'b00000000000000000000101110111100; // input=0.091796875, output=0.091668005704
			11'd24: out = 32'b00000000000000000000110000111011; // input=0.095703125, output=0.0955570996629
			11'd25: out = 32'b00000000000000000000110010111011; // input=0.099609375, output=0.099444735538
			11'd26: out = 32'b00000000000000000000110100111010; // input=0.103515625, output=0.103330854009
			11'd27: out = 32'b00000000000000000000110110111001; // input=0.107421875, output=0.107215395778
			11'd28: out = 32'b00000000000000000000111000111000; // input=0.111328125, output=0.111098301572
			11'd29: out = 32'b00000000000000000000111010111000; // input=0.115234375, output=0.114979512142
			11'd30: out = 32'b00000000000000000000111100110111; // input=0.119140625, output=0.118858968267
			11'd31: out = 32'b00000000000000000000111110110110; // input=0.123046875, output=0.12273661075
			11'd32: out = 32'b00000000000000000001000000110101; // input=0.126953125, output=0.126612380424
			11'd33: out = 32'b00000000000000000001000010110100; // input=0.130859375, output=0.130486218148
			11'd34: out = 32'b00000000000000000001000100110011; // input=0.134765625, output=0.134358064813
			11'd35: out = 32'b00000000000000000001000110110001; // input=0.138671875, output=0.13822786134
			11'd36: out = 32'b00000000000000000001001000110000; // input=0.142578125, output=0.142095548679
			11'd37: out = 32'b00000000000000000001001010101111; // input=0.146484375, output=0.145961067815
			11'd38: out = 32'b00000000000000000001001100101101; // input=0.150390625, output=0.149824359765
			11'd39: out = 32'b00000000000000000001001110101100; // input=0.154296875, output=0.153685365579
			11'd40: out = 32'b00000000000000000001010000101010; // input=0.158203125, output=0.157544026344
			11'd41: out = 32'b00000000000000000001010010101001; // input=0.162109375, output=0.161400283181
			11'd42: out = 32'b00000000000000000001010100100111; // input=0.166015625, output=0.165254077248
			11'd43: out = 32'b00000000000000000001010110100101; // input=0.169921875, output=0.169105349741
			11'd44: out = 32'b00000000000000000001011000100011; // input=0.173828125, output=0.172954041894
			11'd45: out = 32'b00000000000000000001011010100001; // input=0.177734375, output=0.176800094982
			11'd46: out = 32'b00000000000000000001011100011111; // input=0.181640625, output=0.180643450318
			11'd47: out = 32'b00000000000000000001011110011101; // input=0.185546875, output=0.184484049257
			11'd48: out = 32'b00000000000000000001100000011011; // input=0.189453125, output=0.188321833196
			11'd49: out = 32'b00000000000000000001100010011001; // input=0.193359375, output=0.192156743576
			11'd50: out = 32'b00000000000000000001100100010110; // input=0.197265625, output=0.19598872188
			11'd51: out = 32'b00000000000000000001100110010100; // input=0.201171875, output=0.199817709638
			11'd52: out = 32'b00000000000000000001101000010001; // input=0.205078125, output=0.203643648423
			11'd53: out = 32'b00000000000000000001101010001110; // input=0.208984375, output=0.207466479857
			11'd54: out = 32'b00000000000000000001101100001011; // input=0.212890625, output=0.211286145607
			11'd55: out = 32'b00000000000000000001101110001000; // input=0.216796875, output=0.215102587391
			11'd56: out = 32'b00000000000000000001110000000101; // input=0.220703125, output=0.218915746974
			11'd57: out = 32'b00000000000000000001110010000010; // input=0.224609375, output=0.222725566172
			11'd58: out = 32'b00000000000000000001110011111111; // input=0.228515625, output=0.226531986852
			11'd59: out = 32'b00000000000000000001110101111100; // input=0.232421875, output=0.230334950932
			11'd60: out = 32'b00000000000000000001110111111000; // input=0.236328125, output=0.234134400385
			11'd61: out = 32'b00000000000000000001111001110100; // input=0.240234375, output=0.237930277234
			11'd62: out = 32'b00000000000000000001111011110001; // input=0.244140625, output=0.241722523561
			11'd63: out = 32'b00000000000000000001111101101101; // input=0.248046875, output=0.245511081499
			11'd64: out = 32'b00000000000000000001111111101001; // input=0.251953125, output=0.24929589324
			11'd65: out = 32'b00000000000000000010000001100101; // input=0.255859375, output=0.253076901032
			11'd66: out = 32'b00000000000000000010000011100001; // input=0.259765625, output=0.256854047182
			11'd67: out = 32'b00000000000000000010000101011100; // input=0.263671875, output=0.260627274056
			11'd68: out = 32'b00000000000000000010000111011000; // input=0.267578125, output=0.264396524078
			11'd69: out = 32'b00000000000000000010001001010011; // input=0.271484375, output=0.268161739734
			11'd70: out = 32'b00000000000000000010001011001110; // input=0.275390625, output=0.271922863572
			11'd71: out = 32'b00000000000000000010001101001001; // input=0.279296875, output=0.275679838202
			11'd72: out = 32'b00000000000000000010001111000100; // input=0.283203125, output=0.279432606296
			11'd73: out = 32'b00000000000000000010010000111111; // input=0.287109375, output=0.283181110593
			11'd74: out = 32'b00000000000000000010010010111010; // input=0.291015625, output=0.286925293895
			11'd75: out = 32'b00000000000000000010010100110101; // input=0.294921875, output=0.290665099069
			11'd76: out = 32'b00000000000000000010010110101111; // input=0.298828125, output=0.294400469052
			11'd77: out = 32'b00000000000000000010011000101001; // input=0.302734375, output=0.298131346846
			11'd78: out = 32'b00000000000000000010011010100011; // input=0.306640625, output=0.301857675522
			11'd79: out = 32'b00000000000000000010011100011101; // input=0.310546875, output=0.305579398221
			11'd80: out = 32'b00000000000000000010011110010111; // input=0.314453125, output=0.309296458155
			11'd81: out = 32'b00000000000000000010100000010001; // input=0.318359375, output=0.313008798605
			11'd82: out = 32'b00000000000000000010100010001010; // input=0.322265625, output=0.316716362927
			11'd83: out = 32'b00000000000000000010100100000011; // input=0.326171875, output=0.320419094546
			11'd84: out = 32'b00000000000000000010100101111101; // input=0.330078125, output=0.324116936964
			11'd85: out = 32'b00000000000000000010100111110110; // input=0.333984375, output=0.327809833756
			11'd86: out = 32'b00000000000000000010101001101111; // input=0.337890625, output=0.331497728574
			11'd87: out = 32'b00000000000000000010101011100111; // input=0.341796875, output=0.335180565144
			11'd88: out = 32'b00000000000000000010101101100000; // input=0.345703125, output=0.338858287271
			11'd89: out = 32'b00000000000000000010101111011000; // input=0.349609375, output=0.342530838838
			11'd90: out = 32'b00000000000000000010110001010000; // input=0.353515625, output=0.346198163805
			11'd91: out = 32'b00000000000000000010110011001000; // input=0.357421875, output=0.349860206215
			11'd92: out = 32'b00000000000000000010110101000000; // input=0.361328125, output=0.353516910188
			11'd93: out = 32'b00000000000000000010110110111000; // input=0.365234375, output=0.357168219928
			11'd94: out = 32'b00000000000000000010111000101111; // input=0.369140625, output=0.36081407972
			11'd95: out = 32'b00000000000000000010111010100110; // input=0.373046875, output=0.364454433933
			11'd96: out = 32'b00000000000000000010111100011110; // input=0.376953125, output=0.36808922702
			11'd97: out = 32'b00000000000000000010111110010100; // input=0.380859375, output=0.371718403519
			11'd98: out = 32'b00000000000000000011000000001011; // input=0.384765625, output=0.375341908052
			11'd99: out = 32'b00000000000000000011000010000010; // input=0.388671875, output=0.378959685329
			11'd100: out = 32'b00000000000000000011000011111000; // input=0.392578125, output=0.382571680148
			11'd101: out = 32'b00000000000000000011000101101110; // input=0.396484375, output=0.386177837393
			11'd102: out = 32'b00000000000000000011000111100100; // input=0.400390625, output=0.38977810204
			11'd103: out = 32'b00000000000000000011001001011010; // input=0.404296875, output=0.393372419153
			11'd104: out = 32'b00000000000000000011001011010000; // input=0.408203125, output=0.396960733886
			11'd105: out = 32'b00000000000000000011001101000101; // input=0.412109375, output=0.400542991487
			11'd106: out = 32'b00000000000000000011001110111010; // input=0.416015625, output=0.404119137295
			11'd107: out = 32'b00000000000000000011010000101111; // input=0.419921875, output=0.407689116742
			11'd108: out = 32'b00000000000000000011010010100100; // input=0.423828125, output=0.411252875354
			11'd109: out = 32'b00000000000000000011010100011001; // input=0.427734375, output=0.414810358754
			11'd110: out = 32'b00000000000000000011010110001101; // input=0.431640625, output=0.418361512658
			11'd111: out = 32'b00000000000000000011011000000001; // input=0.435546875, output=0.42190628288
			11'd112: out = 32'b00000000000000000011011001110101; // input=0.439453125, output=0.425444615332
			11'd113: out = 32'b00000000000000000011011011101001; // input=0.443359375, output=0.428976456021
			11'd114: out = 32'b00000000000000000011011101011100; // input=0.447265625, output=0.432501751058
			11'd115: out = 32'b00000000000000000011011111010000; // input=0.451171875, output=0.436020446651
			11'd116: out = 32'b00000000000000000011100001000011; // input=0.455078125, output=0.439532489107
			11'd117: out = 32'b00000000000000000011100010110101; // input=0.458984375, output=0.443037824839
			11'd118: out = 32'b00000000000000000011100100101000; // input=0.462890625, output=0.446536400359
			11'd119: out = 32'b00000000000000000011100110011011; // input=0.466796875, output=0.450028162283
			11'd120: out = 32'b00000000000000000011101000001101; // input=0.470703125, output=0.45351305733
			11'd121: out = 32'b00000000000000000011101001111111; // input=0.474609375, output=0.456991032326
			11'd122: out = 32'b00000000000000000011101011110000; // input=0.478515625, output=0.460462034202
			11'd123: out = 32'b00000000000000000011101101100010; // input=0.482421875, output=0.463926009993
			11'd124: out = 32'b00000000000000000011101111010011; // input=0.486328125, output=0.467382906844
			11'd125: out = 32'b00000000000000000011110001000100; // input=0.490234375, output=0.470832672007
			11'd126: out = 32'b00000000000000000011110010110101; // input=0.494140625, output=0.474275252843
			11'd127: out = 32'b00000000000000000011110100100110; // input=0.498046875, output=0.477710596821
			11'd128: out = 32'b00000000000000000011110110010110; // input=0.501953125, output=0.481138651524
			11'd129: out = 32'b00000000000000000011111000000110; // input=0.505859375, output=0.484559364643
			11'd130: out = 32'b00000000000000000011111001110110; // input=0.509765625, output=0.487972683983
			11'd131: out = 32'b00000000000000000011111011100101; // input=0.513671875, output=0.491378557459
			11'd132: out = 32'b00000000000000000011111101010101; // input=0.517578125, output=0.494776933103
			11'd133: out = 32'b00000000000000000011111111000100; // input=0.521484375, output=0.49816775906
			11'd134: out = 32'b00000000000000000100000000110011; // input=0.525390625, output=0.50155098359
			11'd135: out = 32'b00000000000000000100000010100001; // input=0.529296875, output=0.504926555069
			11'd136: out = 32'b00000000000000000100000100010000; // input=0.533203125, output=0.50829442199
			11'd137: out = 32'b00000000000000000100000101111110; // input=0.537109375, output=0.511654532964
			11'd138: out = 32'b00000000000000000100000111101100; // input=0.541015625, output=0.515006836719
			11'd139: out = 32'b00000000000000000100001001011001; // input=0.544921875, output=0.518351282103
			11'd140: out = 32'b00000000000000000100001011000111; // input=0.548828125, output=0.521687818084
			11'd141: out = 32'b00000000000000000100001100110100; // input=0.552734375, output=0.525016393751
			11'd142: out = 32'b00000000000000000100001110100001; // input=0.556640625, output=0.528336958314
			11'd143: out = 32'b00000000000000000100010000001101; // input=0.560546875, output=0.531649461105
			11'd144: out = 32'b00000000000000000100010001111001; // input=0.564453125, output=0.534953851579
			11'd145: out = 32'b00000000000000000100010011100101; // input=0.568359375, output=0.538250079316
			11'd146: out = 32'b00000000000000000100010101010001; // input=0.572265625, output=0.541538094019
			11'd147: out = 32'b00000000000000000100010110111101; // input=0.576171875, output=0.544817845516
			11'd148: out = 32'b00000000000000000100011000101000; // input=0.580078125, output=0.548089283764
			11'd149: out = 32'b00000000000000000100011010010011; // input=0.583984375, output=0.551352358843
			11'd150: out = 32'b00000000000000000100011011111101; // input=0.587890625, output=0.554607020964
			11'd151: out = 32'b00000000000000000100011101101000; // input=0.591796875, output=0.557853220464
			11'd152: out = 32'b00000000000000000100011111010010; // input=0.595703125, output=0.561090907811
			11'd153: out = 32'b00000000000000000100100000111100; // input=0.599609375, output=0.5643200336
			11'd154: out = 32'b00000000000000000100100010100101; // input=0.603515625, output=0.56754054856
			11'd155: out = 32'b00000000000000000100100100001110; // input=0.607421875, output=0.570752403549
			11'd156: out = 32'b00000000000000000100100101110111; // input=0.611328125, output=0.573955549559
			11'd157: out = 32'b00000000000000000100100111100000; // input=0.615234375, output=0.577149937714
			11'd158: out = 32'b00000000000000000100101001001000; // input=0.619140625, output=0.58033551927
			11'd159: out = 32'b00000000000000000100101010110001; // input=0.623046875, output=0.583512245621
			11'd160: out = 32'b00000000000000000100101100011000; // input=0.626953125, output=0.586680068292
			11'd161: out = 32'b00000000000000000100101110000000; // input=0.630859375, output=0.589838938948
			11'd162: out = 32'b00000000000000000100101111100111; // input=0.634765625, output=0.592988809387
			11'd163: out = 32'b00000000000000000100110001001110; // input=0.638671875, output=0.596129631546
			11'd164: out = 32'b00000000000000000100110010110101; // input=0.642578125, output=0.599261357501
			11'd165: out = 32'b00000000000000000100110100011011; // input=0.646484375, output=0.602383939464
			11'd166: out = 32'b00000000000000000100110110000001; // input=0.650390625, output=0.60549732979
			11'd167: out = 32'b00000000000000000100110111100111; // input=0.654296875, output=0.608601480971
			11'd168: out = 32'b00000000000000000100111001001100; // input=0.658203125, output=0.611696345643
			11'd169: out = 32'b00000000000000000100111010110001; // input=0.662109375, output=0.614781876581
			11'd170: out = 32'b00000000000000000100111100010110; // input=0.666015625, output=0.617858026704
			11'd171: out = 32'b00000000000000000100111101111010; // input=0.669921875, output=0.620924749074
			11'd172: out = 32'b00000000000000000100111111011111; // input=0.673828125, output=0.623981996896
			11'd173: out = 32'b00000000000000000101000001000011; // input=0.677734375, output=0.62702972352
			11'd174: out = 32'b00000000000000000101000010100110; // input=0.681640625, output=0.630067882443
			11'd175: out = 32'b00000000000000000101000100001001; // input=0.685546875, output=0.633096427304
			11'd176: out = 32'b00000000000000000101000101101100; // input=0.689453125, output=0.636115311893
			11'd177: out = 32'b00000000000000000101000111001111; // input=0.693359375, output=0.639124490145
			11'd178: out = 32'b00000000000000000101001000110001; // input=0.697265625, output=0.642123916144
			11'd179: out = 32'b00000000000000000101001010010011; // input=0.701171875, output=0.645113544122
			11'd180: out = 32'b00000000000000000101001011110101; // input=0.705078125, output=0.64809332846
			11'd181: out = 32'b00000000000000000101001101010110; // input=0.708984375, output=0.651063223692
			11'd182: out = 32'b00000000000000000101001110110111; // input=0.712890625, output=0.6540231845
			11'd183: out = 32'b00000000000000000101010000011000; // input=0.716796875, output=0.65697316572
			11'd184: out = 32'b00000000000000000101010001111000; // input=0.720703125, output=0.659913122336
			11'd185: out = 32'b00000000000000000101010011011000; // input=0.724609375, output=0.662843009491
			11'd186: out = 32'b00000000000000000101010100111000; // input=0.728515625, output=0.665762782477
			11'd187: out = 32'b00000000000000000101010110010111; // input=0.732421875, output=0.668672396741
			11'd188: out = 32'b00000000000000000101010111110110; // input=0.736328125, output=0.671571807888
			11'd189: out = 32'b00000000000000000101011001010101; // input=0.740234375, output=0.674460971675
			11'd190: out = 32'b00000000000000000101011010110011; // input=0.744140625, output=0.677339844018
			11'd191: out = 32'b00000000000000000101011100010001; // input=0.748046875, output=0.680208380988
			11'd192: out = 32'b00000000000000000101011101101111; // input=0.751953125, output=0.683066538814
			11'd193: out = 32'b00000000000000000101011111001100; // input=0.755859375, output=0.685914273886
			11'd194: out = 32'b00000000000000000101100000101001; // input=0.759765625, output=0.68875154275
			11'd195: out = 32'b00000000000000000101100010000110; // input=0.763671875, output=0.691578302113
			11'd196: out = 32'b00000000000000000101100011100010; // input=0.767578125, output=0.694394508842
			11'd197: out = 32'b00000000000000000101100100111110; // input=0.771484375, output=0.697200119965
			11'd198: out = 32'b00000000000000000101100110011001; // input=0.775390625, output=0.699995092672
			11'd199: out = 32'b00000000000000000101100111110101; // input=0.779296875, output=0.702779384315
			11'd200: out = 32'b00000000000000000101101001010000; // input=0.783203125, output=0.705552952409
			11'd201: out = 32'b00000000000000000101101010101010; // input=0.787109375, output=0.708315754633
			11'd202: out = 32'b00000000000000000101101100000100; // input=0.791015625, output=0.711067748831
			11'd203: out = 32'b00000000000000000101101101011110; // input=0.794921875, output=0.713808893009
			11'd204: out = 32'b00000000000000000101101110111000; // input=0.798828125, output=0.716539145342
			11'd205: out = 32'b00000000000000000101110000010001; // input=0.802734375, output=0.719258464169
			11'd206: out = 32'b00000000000000000101110001101001; // input=0.806640625, output=0.721966807997
			11'd207: out = 32'b00000000000000000101110011000010; // input=0.810546875, output=0.7246641355
			11'd208: out = 32'b00000000000000000101110100011010; // input=0.814453125, output=0.727350405519
			11'd209: out = 32'b00000000000000000101110101110001; // input=0.818359375, output=0.730025577067
			11'd210: out = 32'b00000000000000000101110111001001; // input=0.822265625, output=0.732689609322
			11'd211: out = 32'b00000000000000000101111000100000; // input=0.826171875, output=0.735342461635
			11'd212: out = 32'b00000000000000000101111001110110; // input=0.830078125, output=0.737984093527
			11'd213: out = 32'b00000000000000000101111011001100; // input=0.833984375, output=0.740614464689
			11'd214: out = 32'b00000000000000000101111100100010; // input=0.837890625, output=0.743233534986
			11'd215: out = 32'b00000000000000000101111101111000; // input=0.841796875, output=0.745841264454
			11'd216: out = 32'b00000000000000000101111111001101; // input=0.845703125, output=0.748437613302
			11'd217: out = 32'b00000000000000000110000000100010; // input=0.849609375, output=0.751022541912
			11'd218: out = 32'b00000000000000000110000001110110; // input=0.853515625, output=0.753596010843
			11'd219: out = 32'b00000000000000000110000011001010; // input=0.857421875, output=0.756157980826
			11'd220: out = 32'b00000000000000000110000100011101; // input=0.861328125, output=0.758708412768
			11'd221: out = 32'b00000000000000000110000101110001; // input=0.865234375, output=0.761247267753
			11'd222: out = 32'b00000000000000000110000111000011; // input=0.869140625, output=0.763774507042
			11'd223: out = 32'b00000000000000000110001000010110; // input=0.873046875, output=0.766290092071
			11'd224: out = 32'b00000000000000000110001001101000; // input=0.876953125, output=0.768793984456
			11'd225: out = 32'b00000000000000000110001010111010; // input=0.880859375, output=0.771286145991
			11'd226: out = 32'b00000000000000000110001100001011; // input=0.884765625, output=0.773766538648
			11'd227: out = 32'b00000000000000000110001101011100; // input=0.888671875, output=0.77623512458
			11'd228: out = 32'b00000000000000000110001110101100; // input=0.892578125, output=0.778691866119
			11'd229: out = 32'b00000000000000000110001111111100; // input=0.896484375, output=0.781136725778
			11'd230: out = 32'b00000000000000000110010001001100; // input=0.900390625, output=0.783569666252
			11'd231: out = 32'b00000000000000000110010010011011; // input=0.904296875, output=0.785990650417
			11'd232: out = 32'b00000000000000000110010011101010; // input=0.908203125, output=0.788399641331
			11'd233: out = 32'b00000000000000000110010100111001; // input=0.912109375, output=0.790796602237
			11'd234: out = 32'b00000000000000000110010110000111; // input=0.916015625, output=0.79318149656
			11'd235: out = 32'b00000000000000000110010111010101; // input=0.919921875, output=0.795554287909
			11'd236: out = 32'b00000000000000000110011000100010; // input=0.923828125, output=0.797914940078
			11'd237: out = 32'b00000000000000000110011001101111; // input=0.927734375, output=0.800263417047
			11'd238: out = 32'b00000000000000000110011010111100; // input=0.931640625, output=0.802599682981
			11'd239: out = 32'b00000000000000000110011100001000; // input=0.935546875, output=0.804923702231
			11'd240: out = 32'b00000000000000000110011101010011; // input=0.939453125, output=0.807235439336
			11'd241: out = 32'b00000000000000000110011110011111; // input=0.943359375, output=0.809534859021
			11'd242: out = 32'b00000000000000000110011111101010; // input=0.947265625, output=0.8118219262
			11'd243: out = 32'b00000000000000000110100000110100; // input=0.951171875, output=0.814096605976
			11'd244: out = 32'b00000000000000000110100001111110; // input=0.955078125, output=0.816358863639
			11'd245: out = 32'b00000000000000000110100011001000; // input=0.958984375, output=0.81860866467
			11'd246: out = 32'b00000000000000000110100100010001; // input=0.962890625, output=0.82084597474
			11'd247: out = 32'b00000000000000000110100101011010; // input=0.966796875, output=0.82307075971
			11'd248: out = 32'b00000000000000000110100110100011; // input=0.970703125, output=0.825282985633
			11'd249: out = 32'b00000000000000000110100111101011; // input=0.974609375, output=0.827482618753
			11'd250: out = 32'b00000000000000000110101000110011; // input=0.978515625, output=0.829669625507
			11'd251: out = 32'b00000000000000000110101001111010; // input=0.982421875, output=0.831843972523
			11'd252: out = 32'b00000000000000000110101011000001; // input=0.986328125, output=0.834005626623
			11'd253: out = 32'b00000000000000000110101100000111; // input=0.990234375, output=0.836154554823
			11'd254: out = 32'b00000000000000000110101101001101; // input=0.994140625, output=0.838290724334
			11'd255: out = 32'b00000000000000000110101110010011; // input=0.998046875, output=0.84041410256
			11'd256: out = 32'b00000000000000000110101111011000; // input=1.001953125, output=0.8425246571
			11'd257: out = 32'b00000000000000000110110000011101; // input=1.005859375, output=0.844622355751
			11'd258: out = 32'b00000000000000000110110001100001; // input=1.009765625, output=0.846707166504
			11'd259: out = 32'b00000000000000000110110010100101; // input=1.013671875, output=0.848779057547
			11'd260: out = 32'b00000000000000000110110011101000; // input=1.017578125, output=0.850837997266
			11'd261: out = 32'b00000000000000000110110100101011; // input=1.021484375, output=0.852883954244
			11'd262: out = 32'b00000000000000000110110101101110; // input=1.025390625, output=0.854916897262
			11'd263: out = 32'b00000000000000000110110110110000; // input=1.029296875, output=0.8569367953
			11'd264: out = 32'b00000000000000000110110111110010; // input=1.033203125, output=0.858943617537
			11'd265: out = 32'b00000000000000000110111000110011; // input=1.037109375, output=0.860937333352
			11'd266: out = 32'b00000000000000000110111001110100; // input=1.041015625, output=0.862917912321
			11'd267: out = 32'b00000000000000000110111010110101; // input=1.044921875, output=0.864885324225
			11'd268: out = 32'b00000000000000000110111011110101; // input=1.048828125, output=0.866839539044
			11'd269: out = 32'b00000000000000000110111100110100; // input=1.052734375, output=0.868780526957
			11'd270: out = 32'b00000000000000000110111101110011; // input=1.056640625, output=0.870708258348
			11'd271: out = 32'b00000000000000000110111110110010; // input=1.060546875, output=0.872622703803
			11'd272: out = 32'b00000000000000000110111111110000; // input=1.064453125, output=0.874523834109
			11'd273: out = 32'b00000000000000000111000000101110; // input=1.068359375, output=0.876411620257
			11'd274: out = 32'b00000000000000000111000001101100; // input=1.072265625, output=0.878286033441
			11'd275: out = 32'b00000000000000000111000010101001; // input=1.076171875, output=0.880147045062
			11'd276: out = 32'b00000000000000000111000011100101; // input=1.080078125, output=0.881994626722
			11'd277: out = 32'b00000000000000000111000100100001; // input=1.083984375, output=0.883828750229
			11'd278: out = 32'b00000000000000000111000101011101; // input=1.087890625, output=0.885649387596
			11'd279: out = 32'b00000000000000000111000110011000; // input=1.091796875, output=0.887456511044
			11'd280: out = 32'b00000000000000000111000111010011; // input=1.095703125, output=0.889250092997
			11'd281: out = 32'b00000000000000000111001000001101; // input=1.099609375, output=0.891030106087
			11'd282: out = 32'b00000000000000000111001001000111; // input=1.103515625, output=0.892796523155
			11'd283: out = 32'b00000000000000000111001010000001; // input=1.107421875, output=0.894549317246
			11'd284: out = 32'b00000000000000000111001010111010; // input=1.111328125, output=0.896288461615
			11'd285: out = 32'b00000000000000000111001011110010; // input=1.115234375, output=0.898013929725
			11'd286: out = 32'b00000000000000000111001100101010; // input=1.119140625, output=0.899725695247
			11'd287: out = 32'b00000000000000000111001101100010; // input=1.123046875, output=0.901423732062
			11'd288: out = 32'b00000000000000000111001110011001; // input=1.126953125, output=0.90310801426
			11'd289: out = 32'b00000000000000000111001111010000; // input=1.130859375, output=0.90477851614
			11'd290: out = 32'b00000000000000000111010000000110; // input=1.134765625, output=0.906435212214
			11'd291: out = 32'b00000000000000000111010000111100; // input=1.138671875, output=0.908078077202
			11'd292: out = 32'b00000000000000000111010001110001; // input=1.142578125, output=0.909707086035
			11'd293: out = 32'b00000000000000000111010010100110; // input=1.146484375, output=0.911322213858
			11'd294: out = 32'b00000000000000000111010011011011; // input=1.150390625, output=0.912923436025
			11'd295: out = 32'b00000000000000000111010100001111; // input=1.154296875, output=0.914510728103
			11'd296: out = 32'b00000000000000000111010101000010; // input=1.158203125, output=0.916084065873
			11'd297: out = 32'b00000000000000000111010101110101; // input=1.162109375, output=0.917643425327
			11'd298: out = 32'b00000000000000000111010110101000; // input=1.166015625, output=0.919188782671
			11'd299: out = 32'b00000000000000000111010111011010; // input=1.169921875, output=0.920720114326
			11'd300: out = 32'b00000000000000000111011000001100; // input=1.173828125, output=0.922237396924
			11'd301: out = 32'b00000000000000000111011000111101; // input=1.177734375, output=0.923740607315
			11'd302: out = 32'b00000000000000000111011001101110; // input=1.181640625, output=0.92522972256
			11'd303: out = 32'b00000000000000000111011010011110; // input=1.185546875, output=0.926704719938
			11'd304: out = 32'b00000000000000000111011011001110; // input=1.189453125, output=0.928165576942
			11'd305: out = 32'b00000000000000000111011011111110; // input=1.193359375, output=0.929612271281
			11'd306: out = 32'b00000000000000000111011100101100; // input=1.197265625, output=0.931044780881
			11'd307: out = 32'b00000000000000000111011101011011; // input=1.201171875, output=0.932463083883
			11'd308: out = 32'b00000000000000000111011110001001; // input=1.205078125, output=0.933867158646
			11'd309: out = 32'b00000000000000000111011110110111; // input=1.208984375, output=0.935256983744
			11'd310: out = 32'b00000000000000000111011111100100; // input=1.212890625, output=0.936632537972
			11'd311: out = 32'b00000000000000000111100000010000; // input=1.216796875, output=0.93799380034
			11'd312: out = 32'b00000000000000000111100000111100; // input=1.220703125, output=0.939340750076
			11'd313: out = 32'b00000000000000000111100001101000; // input=1.224609375, output=0.940673366629
			11'd314: out = 32'b00000000000000000111100010010011; // input=1.228515625, output=0.941991629663
			11'd315: out = 32'b00000000000000000111100010111110; // input=1.232421875, output=0.943295519063
			11'd316: out = 32'b00000000000000000111100011101000; // input=1.236328125, output=0.944585014935
			11'd317: out = 32'b00000000000000000111100100010010; // input=1.240234375, output=0.945860097601
			11'd318: out = 32'b00000000000000000111100100111011; // input=1.244140625, output=0.947120747606
			11'd319: out = 32'b00000000000000000111100101100100; // input=1.248046875, output=0.948366945714
			11'd320: out = 32'b00000000000000000111100110001100; // input=1.251953125, output=0.949598672909
			11'd321: out = 32'b00000000000000000111100110110100; // input=1.255859375, output=0.950815910397
			11'd322: out = 32'b00000000000000000111100111011100; // input=1.259765625, output=0.952018639603
			11'd323: out = 32'b00000000000000000111101000000011; // input=1.263671875, output=0.953206842177
			11'd324: out = 32'b00000000000000000111101000101001; // input=1.267578125, output=0.954380499987
			11'd325: out = 32'b00000000000000000111101001001111; // input=1.271484375, output=0.955539595124
			11'd326: out = 32'b00000000000000000111101001110101; // input=1.275390625, output=0.956684109903
			11'd327: out = 32'b00000000000000000111101010011010; // input=1.279296875, output=0.95781402686
			11'd328: out = 32'b00000000000000000111101010111110; // input=1.283203125, output=0.958929328753
			11'd329: out = 32'b00000000000000000111101011100010; // input=1.287109375, output=0.960029998564
			11'd330: out = 32'b00000000000000000111101100000110; // input=1.291015625, output=0.961116019499
			11'd331: out = 32'b00000000000000000111101100101001; // input=1.294921875, output=0.962187374985
			11'd332: out = 32'b00000000000000000111101101001100; // input=1.298828125, output=0.963244048676
			11'd333: out = 32'b00000000000000000111101101101110; // input=1.302734375, output=0.964286024448
			11'd334: out = 32'b00000000000000000111101110001111; // input=1.306640625, output=0.965313286402
			11'd335: out = 32'b00000000000000000111101110110001; // input=1.310546875, output=0.966325818863
			11'd336: out = 32'b00000000000000000111101111010001; // input=1.314453125, output=0.96732360638
			11'd337: out = 32'b00000000000000000111101111110001; // input=1.318359375, output=0.96830663373
			11'd338: out = 32'b00000000000000000111110000010001; // input=1.322265625, output=0.969274885911
			11'd339: out = 32'b00000000000000000111110000110000; // input=1.326171875, output=0.970228348151
			11'd340: out = 32'b00000000000000000111110001001111; // input=1.330078125, output=0.971167005899
			11'd341: out = 32'b00000000000000000111110001101101; // input=1.333984375, output=0.972090844834
			11'd342: out = 32'b00000000000000000111110010001011; // input=1.337890625, output=0.972999850858
			11'd343: out = 32'b00000000000000000111110010101001; // input=1.341796875, output=0.973894010102
			11'd344: out = 32'b00000000000000000111110011000101; // input=1.345703125, output=0.974773308922
			11'd345: out = 32'b00000000000000000111110011100010; // input=1.349609375, output=0.9756377339
			11'd346: out = 32'b00000000000000000111110011111110; // input=1.353515625, output=0.976487271847
			11'd347: out = 32'b00000000000000000111110100011001; // input=1.357421875, output=0.977321909799
			11'd348: out = 32'b00000000000000000111110100110100; // input=1.361328125, output=0.978141635021
			11'd349: out = 32'b00000000000000000111110101001110; // input=1.365234375, output=0.978946435006
			11'd350: out = 32'b00000000000000000111110101101000; // input=1.369140625, output=0.979736297472
			11'd351: out = 32'b00000000000000000111110110000001; // input=1.373046875, output=0.980511210368
			11'd352: out = 32'b00000000000000000111110110011010; // input=1.376953125, output=0.981271161869
			11'd353: out = 32'b00000000000000000111110110110011; // input=1.380859375, output=0.98201614038
			11'd354: out = 32'b00000000000000000111110111001011; // input=1.384765625, output=0.982746134532
			11'd355: out = 32'b00000000000000000111110111100010; // input=1.388671875, output=0.983461133188
			11'd356: out = 32'b00000000000000000111110111111001; // input=1.392578125, output=0.984161125436
			11'd357: out = 32'b00000000000000000111111000001111; // input=1.396484375, output=0.984846100597
			11'd358: out = 32'b00000000000000000111111000100101; // input=1.400390625, output=0.985516048218
			11'd359: out = 32'b00000000000000000111111000111011; // input=1.404296875, output=0.986170958077
			11'd360: out = 32'b00000000000000000111111001010000; // input=1.408203125, output=0.98681082018
			11'd361: out = 32'b00000000000000000111111001100100; // input=1.412109375, output=0.987435624764
			11'd362: out = 32'b00000000000000000111111001111000; // input=1.416015625, output=0.988045362295
			11'd363: out = 32'b00000000000000000111111010001100; // input=1.419921875, output=0.98864002347
			11'd364: out = 32'b00000000000000000111111010011111; // input=1.423828125, output=0.989219599214
			11'd365: out = 32'b00000000000000000111111010110001; // input=1.427734375, output=0.989784080684
			11'd366: out = 32'b00000000000000000111111011000011; // input=1.431640625, output=0.990333459267
			11'd367: out = 32'b00000000000000000111111011010101; // input=1.435546875, output=0.99086772658
			11'd368: out = 32'b00000000000000000111111011100110; // input=1.439453125, output=0.991386874471
			11'd369: out = 32'b00000000000000000111111011110110; // input=1.443359375, output=0.991890895017
			11'd370: out = 32'b00000000000000000111111100000110; // input=1.447265625, output=0.992379780529
			11'd371: out = 32'b00000000000000000111111100010110; // input=1.451171875, output=0.992853523546
			11'd372: out = 32'b00000000000000000111111100100101; // input=1.455078125, output=0.99331211684
			11'd373: out = 32'b00000000000000000111111100110011; // input=1.458984375, output=0.993755553414
			11'd374: out = 32'b00000000000000000111111101000001; // input=1.462890625, output=0.9941838265
			11'd375: out = 32'b00000000000000000111111101001111; // input=1.466796875, output=0.994596929564
			11'd376: out = 32'b00000000000000000111111101011100; // input=1.470703125, output=0.994994856303
			11'd377: out = 32'b00000000000000000111111101101001; // input=1.474609375, output=0.995377600644
			11'd378: out = 32'b00000000000000000111111101110101; // input=1.478515625, output=0.995745156748
			11'd379: out = 32'b00000000000000000111111110000000; // input=1.482421875, output=0.996097519006
			11'd380: out = 32'b00000000000000000111111110001011; // input=1.486328125, output=0.996434682041
			11'd381: out = 32'b00000000000000000111111110010110; // input=1.490234375, output=0.996756640709
			11'd382: out = 32'b00000000000000000111111110100000; // input=1.494140625, output=0.997063390097
			11'd383: out = 32'b00000000000000000111111110101001; // input=1.498046875, output=0.997354925525
			11'd384: out = 32'b00000000000000000111111110110010; // input=1.501953125, output=0.997631242543
			11'd385: out = 32'b00000000000000000111111110111011; // input=1.505859375, output=0.997892336936
			11'd386: out = 32'b00000000000000000111111111000011; // input=1.509765625, output=0.99813820472
			11'd387: out = 32'b00000000000000000111111111001011; // input=1.513671875, output=0.998368842143
			11'd388: out = 32'b00000000000000000111111111010010; // input=1.517578125, output=0.998584245685
			11'd389: out = 32'b00000000000000000111111111011000; // input=1.521484375, output=0.998784412061
			11'd390: out = 32'b00000000000000000111111111011110; // input=1.525390625, output=0.998969338215
			11'd391: out = 32'b00000000000000000111111111100100; // input=1.529296875, output=0.999139021326
			11'd392: out = 32'b00000000000000000111111111101001; // input=1.533203125, output=0.999293458805
			11'd393: out = 32'b00000000000000000111111111101101; // input=1.537109375, output=0.999432648295
			11'd394: out = 32'b00000000000000000111111111110001; // input=1.541015625, output=0.999556587673
			11'd395: out = 32'b00000000000000000111111111110101; // input=1.544921875, output=0.999665275047
			11'd396: out = 32'b00000000000000000111111111111000; // input=1.548828125, output=0.999758708759
			11'd397: out = 32'b00000000000000000111111111111011; // input=1.552734375, output=0.999836887383
			11'd398: out = 32'b00000000000000000111111111111101; // input=1.556640625, output=0.999899809726
			11'd399: out = 32'b00000000000000000111111111111110; // input=1.560546875, output=0.999947474829
			11'd400: out = 32'b00000000000000000111111111111111; // input=1.564453125, output=0.999979881963
			11'd401: out = 32'b00000000000000000111111111111111; // input=1.568359375, output=0.999997030634
			11'd402: out = 32'b00000000000000000111111111111111; // input=1.572265625, output=0.999998920582
			11'd403: out = 32'b00000000000000000111111111111111; // input=1.576171875, output=0.999985551776
			11'd404: out = 32'b00000000000000000111111111111111; // input=1.580078125, output=0.99995692442
			11'd405: out = 32'b00000000000000000111111111111101; // input=1.583984375, output=0.999913038953
			11'd406: out = 32'b00000000000000000111111111111011; // input=1.587890625, output=0.999853896042
			11'd407: out = 32'b00000000000000000111111111111001; // input=1.591796875, output=0.999779496592
			11'd408: out = 32'b00000000000000000111111111110110; // input=1.595703125, output=0.999689841736
			11'd409: out = 32'b00000000000000000111111111110010; // input=1.599609375, output=0.999584932843
			11'd410: out = 32'b00000000000000000111111111101110; // input=1.603515625, output=0.999464771514
			11'd411: out = 32'b00000000000000000111111111101010; // input=1.607421875, output=0.999329359583
			11'd412: out = 32'b00000000000000000111111111100101; // input=1.611328125, output=0.999178699114
			11'd413: out = 32'b00000000000000000111111111100000; // input=1.615234375, output=0.999012792408
			11'd414: out = 32'b00000000000000000111111111011010; // input=1.619140625, output=0.998831641997
			11'd415: out = 32'b00000000000000000111111111010011; // input=1.623046875, output=0.998635250643
			11'd416: out = 32'b00000000000000000111111111001100; // input=1.626953125, output=0.998423621343
			11'd417: out = 32'b00000000000000000111111111000101; // input=1.630859375, output=0.998196757328
			11'd418: out = 32'b00000000000000000111111110111101; // input=1.634765625, output=0.997954662059
			11'd419: out = 32'b00000000000000000111111110110101; // input=1.638671875, output=0.997697339229
			11'd420: out = 32'b00000000000000000111111110101100; // input=1.642578125, output=0.997424792765
			11'd421: out = 32'b00000000000000000111111110100010; // input=1.646484375, output=0.997137026826
			11'd422: out = 32'b00000000000000000111111110011000; // input=1.650390625, output=0.996834045803
			11'd423: out = 32'b00000000000000000111111110001110; // input=1.654296875, output=0.996515854318
			11'd424: out = 32'b00000000000000000111111110000011; // input=1.658203125, output=0.996182457228
			11'd425: out = 32'b00000000000000000111111101110111; // input=1.662109375, output=0.995833859619
			11'd426: out = 32'b00000000000000000111111101101100; // input=1.666015625, output=0.995470066811
			11'd427: out = 32'b00000000000000000111111101011111; // input=1.669921875, output=0.995091084354
			11'd428: out = 32'b00000000000000000111111101010010; // input=1.673828125, output=0.994696918032
			11'd429: out = 32'b00000000000000000111111101000101; // input=1.677734375, output=0.994287573858
			11'd430: out = 32'b00000000000000000111111100110111; // input=1.681640625, output=0.99386305808
			11'd431: out = 32'b00000000000000000111111100101000; // input=1.685546875, output=0.993423377174
			11'd432: out = 32'b00000000000000000111111100011010; // input=1.689453125, output=0.992968537849
			11'd433: out = 32'b00000000000000000111111100001010; // input=1.693359375, output=0.992498547046
			11'd434: out = 32'b00000000000000000111111011111010; // input=1.697265625, output=0.992013411937
			11'd435: out = 32'b00000000000000000111111011101010; // input=1.701171875, output=0.991513139923
			11'd436: out = 32'b00000000000000000111111011011001; // input=1.705078125, output=0.990997738639
			11'd437: out = 32'b00000000000000000111111011001000; // input=1.708984375, output=0.990467215948
			11'd438: out = 32'b00000000000000000111111010110110; // input=1.712890625, output=0.989921579947
			11'd439: out = 32'b00000000000000000111111010100011; // input=1.716796875, output=0.98936083896
			11'd440: out = 32'b00000000000000000111111010010001; // input=1.720703125, output=0.988785001544
			11'd441: out = 32'b00000000000000000111111001111101; // input=1.724609375, output=0.988194076485
			11'd442: out = 32'b00000000000000000111111001101001; // input=1.728515625, output=0.9875880728
			11'd443: out = 32'b00000000000000000111111001010101; // input=1.732421875, output=0.986966999737
			11'd444: out = 32'b00000000000000000111111001000000; // input=1.736328125, output=0.986330866772
			11'd445: out = 32'b00000000000000000111111000101011; // input=1.740234375, output=0.98567968361
			11'd446: out = 32'b00000000000000000111111000010101; // input=1.744140625, output=0.98501346019
			11'd447: out = 32'b00000000000000000111110111111111; // input=1.748046875, output=0.984332206676
			11'd448: out = 32'b00000000000000000111110111101000; // input=1.751953125, output=0.983635933464
			11'd449: out = 32'b00000000000000000111110111010000; // input=1.755859375, output=0.982924651178
			11'd450: out = 32'b00000000000000000111110110111001; // input=1.759765625, output=0.982198370671
			11'd451: out = 32'b00000000000000000111110110100000; // input=1.763671875, output=0.981457103025
			11'd452: out = 32'b00000000000000000111110110001000; // input=1.767578125, output=0.980700859551
			11'd453: out = 32'b00000000000000000111110101101110; // input=1.771484375, output=0.979929651789
			11'd454: out = 32'b00000000000000000111110101010101; // input=1.775390625, output=0.979143491506
			11'd455: out = 32'b00000000000000000111110100111010; // input=1.779296875, output=0.978342390698
			11'd456: out = 32'b00000000000000000111110100100000; // input=1.783203125, output=0.977526361588
			11'd457: out = 32'b00000000000000000111110100000100; // input=1.787109375, output=0.976695416629
			11'd458: out = 32'b00000000000000000111110011101001; // input=1.791015625, output=0.9758495685
			11'd459: out = 32'b00000000000000000111110011001100; // input=1.794921875, output=0.974988830107
			11'd460: out = 32'b00000000000000000111110010110000; // input=1.798828125, output=0.974113214584
			11'd461: out = 32'b00000000000000000111110010010011; // input=1.802734375, output=0.973222735292
			11'd462: out = 32'b00000000000000000111110001110101; // input=1.806640625, output=0.972317405818
			11'd463: out = 32'b00000000000000000111110001010111; // input=1.810546875, output=0.971397239977
			11'd464: out = 32'b00000000000000000111110000111000; // input=1.814453125, output=0.970462251809
			11'd465: out = 32'b00000000000000000111110000011001; // input=1.818359375, output=0.969512455581
			11'd466: out = 32'b00000000000000000111101111111001; // input=1.822265625, output=0.968547865786
			11'd467: out = 32'b00000000000000000111101111011001; // input=1.826171875, output=0.967568497142
			11'd468: out = 32'b00000000000000000111101110111001; // input=1.830078125, output=0.966574364594
			11'd469: out = 32'b00000000000000000111101110011000; // input=1.833984375, output=0.96556548331
			11'd470: out = 32'b00000000000000000111101101110110; // input=1.837890625, output=0.964541868684
			11'd471: out = 32'b00000000000000000111101101010100; // input=1.841796875, output=0.963503536336
			11'd472: out = 32'b00000000000000000111101100110010; // input=1.845703125, output=0.96245050211
			11'd473: out = 32'b00000000000000000111101100001111; // input=1.849609375, output=0.961382782073
			11'd474: out = 32'b00000000000000000111101011101011; // input=1.853515625, output=0.960300392518
			11'd475: out = 32'b00000000000000000111101011000111; // input=1.857421875, output=0.95920334996
			11'd476: out = 32'b00000000000000000111101010100011; // input=1.861328125, output=0.95809167114
			11'd477: out = 32'b00000000000000000111101001111110; // input=1.865234375, output=0.956965373019
			11'd478: out = 32'b00000000000000000111101001011000; // input=1.869140625, output=0.955824472784
			11'd479: out = 32'b00000000000000000111101000110011; // input=1.873046875, output=0.954668987843
			11'd480: out = 32'b00000000000000000111101000001100; // input=1.876953125, output=0.953498935829
			11'd481: out = 32'b00000000000000000111100111100101; // input=1.880859375, output=0.952314334593
			11'd482: out = 32'b00000000000000000111100110111110; // input=1.884765625, output=0.951115202213
			11'd483: out = 32'b00000000000000000111100110010110; // input=1.888671875, output=0.949901556985
			11'd484: out = 32'b00000000000000000111100101101110; // input=1.892578125, output=0.948673417428
			11'd485: out = 32'b00000000000000000111100101000101; // input=1.896484375, output=0.947430802281
			11'd486: out = 32'b00000000000000000111100100011100; // input=1.900390625, output=0.946173730507
			11'd487: out = 32'b00000000000000000111100011110011; // input=1.904296875, output=0.944902221285
			11'd488: out = 32'b00000000000000000111100011001000; // input=1.908203125, output=0.943616294018
			11'd489: out = 32'b00000000000000000111100010011110; // input=1.912109375, output=0.942315968327
			11'd490: out = 32'b00000000000000000111100001110011; // input=1.916015625, output=0.941001264054
			11'd491: out = 32'b00000000000000000111100001000111; // input=1.919921875, output=0.939672201259
			11'd492: out = 32'b00000000000000000111100000011011; // input=1.923828125, output=0.938328800223
			11'd493: out = 32'b00000000000000000111011111101111; // input=1.927734375, output=0.936971081444
			11'd494: out = 32'b00000000000000000111011111000010; // input=1.931640625, output=0.935599065638
			11'd495: out = 32'b00000000000000000111011110010100; // input=1.935546875, output=0.934212773742
			11'd496: out = 32'b00000000000000000111011101100110; // input=1.939453125, output=0.932812226909
			11'd497: out = 32'b00000000000000000111011100111000; // input=1.943359375, output=0.931397446509
			11'd498: out = 32'b00000000000000000111011100001001; // input=1.947265625, output=0.929968454129
			11'd499: out = 32'b00000000000000000111011011011010; // input=1.951171875, output=0.928525271575
			11'd500: out = 32'b00000000000000000111011010101010; // input=1.955078125, output=0.927067920868
			11'd501: out = 32'b00000000000000000111011001111010; // input=1.958984375, output=0.925596424245
			11'd502: out = 32'b00000000000000000111011001001001; // input=1.962890625, output=0.92411080416
			11'd503: out = 32'b00000000000000000111011000011000; // input=1.966796875, output=0.92261108328
			11'd504: out = 32'b00000000000000000111010111100111; // input=1.970703125, output=0.921097284491
			11'd505: out = 32'b00000000000000000111010110110100; // input=1.974609375, output=0.91956943089
			11'd506: out = 32'b00000000000000000111010110000010; // input=1.978515625, output=0.918027545791
			11'd507: out = 32'b00000000000000000111010101001111; // input=1.982421875, output=0.916471652721
			11'd508: out = 32'b00000000000000000111010100011100; // input=1.986328125, output=0.914901775422
			11'd509: out = 32'b00000000000000000111010011101000; // input=1.990234375, output=0.913317937847
			11'd510: out = 32'b00000000000000000111010010110011; // input=1.994140625, output=0.911720164164
			11'd511: out = 32'b00000000000000000111010001111110; // input=1.998046875, output=0.910108478752
			11'd512: out = 32'b00000000000000000111010001001001; // input=2.001953125, output=0.908482906206
			11'd513: out = 32'b00000000000000000111010000010011; // input=2.005859375, output=0.906843471327
			11'd514: out = 32'b00000000000000000111001111011101; // input=2.009765625, output=0.905190199134
			11'd515: out = 32'b00000000000000000111001110100111; // input=2.013671875, output=0.903523114851
			11'd516: out = 32'b00000000000000000111001101110000; // input=2.017578125, output=0.901842243918
			11'd517: out = 32'b00000000000000000111001100111000; // input=2.021484375, output=0.900147611981
			11'd518: out = 32'b00000000000000000111001100000000; // input=2.025390625, output=0.898439244899
			11'd519: out = 32'b00000000000000000111001011001000; // input=2.029296875, output=0.89671716874
			11'd520: out = 32'b00000000000000000111001010001111; // input=2.033203125, output=0.89498140978
			11'd521: out = 32'b00000000000000000111001001010101; // input=2.037109375, output=0.893231994505
			11'd522: out = 32'b00000000000000000111001000011100; // input=2.041015625, output=0.891468949608
			11'd523: out = 32'b00000000000000000111000111100001; // input=2.044921875, output=0.889692301992
			11'd524: out = 32'b00000000000000000111000110100111; // input=2.048828125, output=0.887902078767
			11'd525: out = 32'b00000000000000000111000101101100; // input=2.052734375, output=0.886098307248
			11'd526: out = 32'b00000000000000000111000100110000; // input=2.056640625, output=0.884281014959
			11'd527: out = 32'b00000000000000000111000011110100; // input=2.060546875, output=0.882450229629
			11'd528: out = 32'b00000000000000000111000010111000; // input=2.064453125, output=0.880605979195
			11'd529: out = 32'b00000000000000000111000001111011; // input=2.068359375, output=0.878748291797
			11'd530: out = 32'b00000000000000000111000000111110; // input=2.072265625, output=0.876877195782
			11'd531: out = 32'b00000000000000000111000000000000; // input=2.076171875, output=0.874992719699
			11'd532: out = 32'b00000000000000000110111111000010; // input=2.080078125, output=0.873094892304
			11'd533: out = 32'b00000000000000000110111110000011; // input=2.083984375, output=0.871183742555
			11'd534: out = 32'b00000000000000000110111101000100; // input=2.087890625, output=0.869259299614
			11'd535: out = 32'b00000000000000000110111100000100; // input=2.091796875, output=0.867321592845
			11'd536: out = 32'b00000000000000000110111011000100; // input=2.095703125, output=0.865370651816
			11'd537: out = 32'b00000000000000000110111010000100; // input=2.099609375, output=0.863406506296
			11'd538: out = 32'b00000000000000000110111001000011; // input=2.103515625, output=0.861429186254
			11'd539: out = 32'b00000000000000000110111000000010; // input=2.107421875, output=0.859438721864
			11'd540: out = 32'b00000000000000000110110111000000; // input=2.111328125, output=0.857435143495
			11'd541: out = 32'b00000000000000000110110101111110; // input=2.115234375, output=0.855418481721
			11'd542: out = 32'b00000000000000000110110100111100; // input=2.119140625, output=0.853388767314
			11'd543: out = 32'b00000000000000000110110011111001; // input=2.123046875, output=0.851346031244
			11'd544: out = 32'b00000000000000000110110010110110; // input=2.126953125, output=0.849290304681
			11'd545: out = 32'b00000000000000000110110001110010; // input=2.130859375, output=0.847221618993
			11'd546: out = 32'b00000000000000000110110000101110; // input=2.134765625, output=0.845140005746
			11'd547: out = 32'b00000000000000000110101111101001; // input=2.138671875, output=0.843045496701
			11'd548: out = 32'b00000000000000000110101110100100; // input=2.142578125, output=0.84093812382
			11'd549: out = 32'b00000000000000000110101101011110; // input=2.146484375, output=0.838817919257
			11'd550: out = 32'b00000000000000000110101100011000; // input=2.150390625, output=0.836684915366
			11'd551: out = 32'b00000000000000000110101011010010; // input=2.154296875, output=0.834539144691
			11'd552: out = 32'b00000000000000000110101010001011; // input=2.158203125, output=0.832380639976
			11'd553: out = 32'b00000000000000000110101001000100; // input=2.162109375, output=0.830209434157
			11'd554: out = 32'b00000000000000000110100111111101; // input=2.166015625, output=0.828025560363
			11'd555: out = 32'b00000000000000000110100110110101; // input=2.169921875, output=0.825829051918
			11'd556: out = 32'b00000000000000000110100101101100; // input=2.173828125, output=0.823619942338
			11'd557: out = 32'b00000000000000000110100100100100; // input=2.177734375, output=0.82139826533
			11'd558: out = 32'b00000000000000000110100011011010; // input=2.181640625, output=0.819164054796
			11'd559: out = 32'b00000000000000000110100010010001; // input=2.185546875, output=0.816917344826
			11'd560: out = 32'b00000000000000000110100001000111; // input=2.189453125, output=0.814658169702
			11'd561: out = 32'b00000000000000000110011111111100; // input=2.193359375, output=0.812386563897
			11'd562: out = 32'b00000000000000000110011110110001; // input=2.197265625, output=0.810102562073
			11'd563: out = 32'b00000000000000000110011101100110; // input=2.201171875, output=0.80780619908
			11'd564: out = 32'b00000000000000000110011100011011; // input=2.205078125, output=0.805497509959
			11'd565: out = 32'b00000000000000000110011011001110; // input=2.208984375, output=0.803176529936
			11'd566: out = 32'b00000000000000000110011010000010; // input=2.212890625, output=0.800843294428
			11'd567: out = 32'b00000000000000000110011000110101; // input=2.216796875, output=0.798497839037
			11'd568: out = 32'b00000000000000000110010111101000; // input=2.220703125, output=0.796140199551
			11'd569: out = 32'b00000000000000000110010110011010; // input=2.224609375, output=0.793770411945
			11'd570: out = 32'b00000000000000000110010101001100; // input=2.228515625, output=0.791388512379
			11'd571: out = 32'b00000000000000000110010011111110; // input=2.232421875, output=0.788994537198
			11'd572: out = 32'b00000000000000000110010010101111; // input=2.236328125, output=0.786588522931
			11'd573: out = 32'b00000000000000000110010001100000; // input=2.240234375, output=0.784170506291
			11'd574: out = 32'b00000000000000000110010000010000; // input=2.244140625, output=0.781740524174
			11'd575: out = 32'b00000000000000000110001111000000; // input=2.248046875, output=0.779298613658
			11'd576: out = 32'b00000000000000000110001101110000; // input=2.251953125, output=0.776844812005
			11'd577: out = 32'b00000000000000000110001100011111; // input=2.255859375, output=0.774379156655
			11'd578: out = 32'b00000000000000000110001011001110; // input=2.259765625, output=0.771901685232
			11'd579: out = 32'b00000000000000000110001001111100; // input=2.263671875, output=0.769412435539
			11'd580: out = 32'b00000000000000000110001000101010; // input=2.267578125, output=0.766911445559
			11'd581: out = 32'b00000000000000000110000111011000; // input=2.271484375, output=0.764398753454
			11'd582: out = 32'b00000000000000000110000110000101; // input=2.275390625, output=0.761874397564
			11'd583: out = 32'b00000000000000000110000100110010; // input=2.279296875, output=0.759338416409
			11'd584: out = 32'b00000000000000000110000011011111; // input=2.283203125, output=0.756790848683
			11'd585: out = 32'b00000000000000000110000010001011; // input=2.287109375, output=0.75423173326
			11'd586: out = 32'b00000000000000000110000000110110; // input=2.291015625, output=0.751661109189
			11'd587: out = 32'b00000000000000000101111111100010; // input=2.294921875, output=0.749079015694
			11'd588: out = 32'b00000000000000000101111110001101; // input=2.298828125, output=0.746485492175
			11'd589: out = 32'b00000000000000000101111100110111; // input=2.302734375, output=0.743880578206
			11'd590: out = 32'b00000000000000000101111011100010; // input=2.306640625, output=0.741264313535
			11'd591: out = 32'b00000000000000000101111010001100; // input=2.310546875, output=0.738636738082
			11'd592: out = 32'b00000000000000000101111000110101; // input=2.314453125, output=0.735997891941
			11'd593: out = 32'b00000000000000000101110111011110; // input=2.318359375, output=0.733347815378
			11'd594: out = 32'b00000000000000000101110110000111; // input=2.322265625, output=0.730686548829
			11'd595: out = 32'b00000000000000000101110100110000; // input=2.326171875, output=0.728014132903
			11'd596: out = 32'b00000000000000000101110011011000; // input=2.330078125, output=0.725330608377
			11'd597: out = 32'b00000000000000000101110001111111; // input=2.333984375, output=0.722636016198
			11'd598: out = 32'b00000000000000000101110000100111; // input=2.337890625, output=0.719930397482
			11'd599: out = 32'b00000000000000000101101111001110; // input=2.341796875, output=0.717213793515
			11'd600: out = 32'b00000000000000000101101101110100; // input=2.345703125, output=0.714486245747
			11'd601: out = 32'b00000000000000000101101100011011; // input=2.349609375, output=0.711747795798
			11'd602: out = 32'b00000000000000000101101011000000; // input=2.353515625, output=0.708998485454
			11'd603: out = 32'b00000000000000000101101001100110; // input=2.357421875, output=0.706238356665
			11'd604: out = 32'b00000000000000000101101000001011; // input=2.361328125, output=0.703467451548
			11'd605: out = 32'b00000000000000000101100110110000; // input=2.365234375, output=0.700685812383
			11'd606: out = 32'b00000000000000000101100101010101; // input=2.369140625, output=0.697893481614
			11'd607: out = 32'b00000000000000000101100011111001; // input=2.373046875, output=0.69509050185
			11'd608: out = 32'b00000000000000000101100010011101; // input=2.376953125, output=0.692276915859
			11'd609: out = 32'b00000000000000000101100001000000; // input=2.380859375, output=0.689452766575
			11'd610: out = 32'b00000000000000000101011111100011; // input=2.384765625, output=0.68661809709
			11'd611: out = 32'b00000000000000000101011110000110; // input=2.388671875, output=0.683772950657
			11'd612: out = 32'b00000000000000000101011100101000; // input=2.392578125, output=0.680917370691
			11'd613: out = 32'b00000000000000000101011011001010; // input=2.396484375, output=0.678051400763
			11'd614: out = 32'b00000000000000000101011001101100; // input=2.400390625, output=0.675175084605
			11'd615: out = 32'b00000000000000000101011000001110; // input=2.404296875, output=0.672288466105
			11'd616: out = 32'b00000000000000000101010110101111; // input=2.408203125, output=0.669391589311
			11'd617: out = 32'b00000000000000000101010101001111; // input=2.412109375, output=0.666484498425
			11'd618: out = 32'b00000000000000000101010011110000; // input=2.416015625, output=0.663567237806
			11'd619: out = 32'b00000000000000000101010010010000; // input=2.419921875, output=0.660639851967
			11'd620: out = 32'b00000000000000000101010000110000; // input=2.423828125, output=0.657702385576
			11'd621: out = 32'b00000000000000000101001111001111; // input=2.427734375, output=0.654754883457
			11'd622: out = 32'b00000000000000000101001101101110; // input=2.431640625, output=0.651797390583
			11'd623: out = 32'b00000000000000000101001100001101; // input=2.435546875, output=0.648829952083
			11'd624: out = 32'b00000000000000000101001010101011; // input=2.439453125, output=0.645852613236
			11'd625: out = 32'b00000000000000000101001001001001; // input=2.443359375, output=0.642865419473
			11'd626: out = 32'b00000000000000000101000111100111; // input=2.447265625, output=0.639868416375
			11'd627: out = 32'b00000000000000000101000110000101; // input=2.451171875, output=0.636861649672
			11'd628: out = 32'b00000000000000000101000100100010; // input=2.455078125, output=0.633845165244
			11'd629: out = 32'b00000000000000000101000010111111; // input=2.458984375, output=0.630819009118
			11'd630: out = 32'b00000000000000000101000001011011; // input=2.462890625, output=0.62778322747
			11'd631: out = 32'b00000000000000000100111111110111; // input=2.466796875, output=0.624737866623
			11'd632: out = 32'b00000000000000000100111110010011; // input=2.470703125, output=0.621682973045
			11'd633: out = 32'b00000000000000000100111100101111; // input=2.474609375, output=0.618618593349
			11'd634: out = 32'b00000000000000000100111011001010; // input=2.478515625, output=0.615544774295
			11'd635: out = 32'b00000000000000000100111001100101; // input=2.482421875, output=0.612461562784
			11'd636: out = 32'b00000000000000000100111000000000; // input=2.486328125, output=0.609369005864
			11'd637: out = 32'b00000000000000000100110110011010; // input=2.490234375, output=0.606267150722
			11'd638: out = 32'b00000000000000000100110100110100; // input=2.494140625, output=0.60315604469
			11'd639: out = 32'b00000000000000000100110011001110; // input=2.498046875, output=0.600035735239
			11'd640: out = 32'b00000000000000000100110001100111; // input=2.501953125, output=0.59690626998
			11'd641: out = 32'b00000000000000000100110000000001; // input=2.505859375, output=0.593767696666
			11'd642: out = 32'b00000000000000000100101110011001; // input=2.509765625, output=0.590620063188
			11'd643: out = 32'b00000000000000000100101100110010; // input=2.513671875, output=0.587463417574
			11'd644: out = 32'b00000000000000000100101011001010; // input=2.517578125, output=0.584297807991
			11'd645: out = 32'b00000000000000000100101001100010; // input=2.521484375, output=0.581123282743
			11'd646: out = 32'b00000000000000000100100111111010; // input=2.525390625, output=0.577939890268
			11'd647: out = 32'b00000000000000000100100110010001; // input=2.529296875, output=0.574747679141
			11'd648: out = 32'b00000000000000000100100100101000; // input=2.533203125, output=0.571546698072
			11'd649: out = 32'b00000000000000000100100010111111; // input=2.537109375, output=0.568336995904
			11'd650: out = 32'b00000000000000000100100001010110; // input=2.541015625, output=0.565118621612
			11'd651: out = 32'b00000000000000000100011111101100; // input=2.544921875, output=0.561891624306
			11'd652: out = 32'b00000000000000000100011110000010; // input=2.548828125, output=0.558656053224
			11'd653: out = 32'b00000000000000000100011100011000; // input=2.552734375, output=0.555411957739
			11'd654: out = 32'b00000000000000000100011010101101; // input=2.556640625, output=0.55215938735
			11'd655: out = 32'b00000000000000000100011001000010; // input=2.560546875, output=0.548898391689
			11'd656: out = 32'b00000000000000000100010111010111; // input=2.564453125, output=0.545629020513
			11'd657: out = 32'b00000000000000000100010101101100; // input=2.568359375, output=0.54235132371
			11'd658: out = 32'b00000000000000000100010100000000; // input=2.572265625, output=0.539065351293
			11'd659: out = 32'b00000000000000000100010010010100; // input=2.576171875, output=0.535771153402
			11'd660: out = 32'b00000000000000000100010000101000; // input=2.580078125, output=0.532468780302
			11'd661: out = 32'b00000000000000000100001110111011; // input=2.583984375, output=0.529158282384
			11'd662: out = 32'b00000000000000000100001101001111; // input=2.587890625, output=0.525839710162
			11'd663: out = 32'b00000000000000000100001011100010; // input=2.591796875, output=0.522513114272
			11'd664: out = 32'b00000000000000000100001001110100; // input=2.595703125, output=0.519178545475
			11'd665: out = 32'b00000000000000000100001000000111; // input=2.599609375, output=0.515836054653
			11'd666: out = 32'b00000000000000000100000110011001; // input=2.603515625, output=0.512485692806
			11'd667: out = 32'b00000000000000000100000100101011; // input=2.607421875, output=0.509127511059
			11'd668: out = 32'b00000000000000000100000010111101; // input=2.611328125, output=0.505761560652
			11'd669: out = 32'b00000000000000000100000001001110; // input=2.615234375, output=0.502387892946
			11'd670: out = 32'b00000000000000000011111111011111; // input=2.619140625, output=0.499006559419
			11'd671: out = 32'b00000000000000000011111101110000; // input=2.623046875, output=0.495617611666
			11'd672: out = 32'b00000000000000000011111100000001; // input=2.626953125, output=0.492221101398
			11'd673: out = 32'b00000000000000000011111010010010; // input=2.630859375, output=0.488817080442
			11'd674: out = 32'b00000000000000000011111000100010; // input=2.634765625, output=0.485405600738
			11'd675: out = 32'b00000000000000000011110110110010; // input=2.638671875, output=0.481986714342
			11'd676: out = 32'b00000000000000000011110101000001; // input=2.642578125, output=0.478560473421
			11'd677: out = 32'b00000000000000000011110011010001; // input=2.646484375, output=0.475126930257
			11'd678: out = 32'b00000000000000000011110001100000; // input=2.650390625, output=0.47168613724
			11'd679: out = 32'b00000000000000000011101111101111; // input=2.654296875, output=0.468238146873
			11'd680: out = 32'b00000000000000000011101101111110; // input=2.658203125, output=0.464783011769
			11'd681: out = 32'b00000000000000000011101100001101; // input=2.662109375, output=0.461320784647
			11'd682: out = 32'b00000000000000000011101010011011; // input=2.666015625, output=0.457851518337
			11'd683: out = 32'b00000000000000000011101000101001; // input=2.669921875, output=0.454375265777
			11'd684: out = 32'b00000000000000000011100110110111; // input=2.673828125, output=0.450892080009
			11'd685: out = 32'b00000000000000000011100101000100; // input=2.677734375, output=0.447402014183
			11'd686: out = 32'b00000000000000000011100011010010; // input=2.681640625, output=0.443905121553
			11'd687: out = 32'b00000000000000000011100001011111; // input=2.685546875, output=0.440401455476
			11'd688: out = 32'b00000000000000000011011111101100; // input=2.689453125, output=0.436891069416
			11'd689: out = 32'b00000000000000000011011101111001; // input=2.693359375, output=0.433374016935
			11'd690: out = 32'b00000000000000000011011100000101; // input=2.697265625, output=0.429850351699
			11'd691: out = 32'b00000000000000000011011010010010; // input=2.701171875, output=0.426320127476
			11'd692: out = 32'b00000000000000000011011000011110; // input=2.705078125, output=0.422783398133
			11'd693: out = 32'b00000000000000000011010110101010; // input=2.708984375, output=0.419240217635
			11'd694: out = 32'b00000000000000000011010100110101; // input=2.712890625, output=0.415690640047
			11'd695: out = 32'b00000000000000000011010011000001; // input=2.716796875, output=0.412134719532
			11'd696: out = 32'b00000000000000000011010001001100; // input=2.720703125, output=0.408572510347
			11'd697: out = 32'b00000000000000000011001111010111; // input=2.724609375, output=0.405004066849
			11'd698: out = 32'b00000000000000000011001101100010; // input=2.728515625, output=0.401429443487
			11'd699: out = 32'b00000000000000000011001011101101; // input=2.732421875, output=0.397848694806
			11'd700: out = 32'b00000000000000000011001001110111; // input=2.736328125, output=0.394261875443
			11'd701: out = 32'b00000000000000000011001000000001; // input=2.740234375, output=0.390669040129
			11'd702: out = 32'b00000000000000000011000110001100; // input=2.744140625, output=0.387070243686
			11'd703: out = 32'b00000000000000000011000100010101; // input=2.748046875, output=0.383465541027
			11'd704: out = 32'b00000000000000000011000010011111; // input=2.751953125, output=0.379854987156
			11'd705: out = 32'b00000000000000000011000000101001; // input=2.755859375, output=0.376238637166
			11'd706: out = 32'b00000000000000000010111110110010; // input=2.759765625, output=0.372616546236
			11'd707: out = 32'b00000000000000000010111100111011; // input=2.763671875, output=0.368988769637
			11'd708: out = 32'b00000000000000000010111011000100; // input=2.767578125, output=0.365355362723
			11'd709: out = 32'b00000000000000000010111001001101; // input=2.771484375, output=0.361716380935
			11'd710: out = 32'b00000000000000000010110111010101; // input=2.775390625, output=0.358071879801
			11'd711: out = 32'b00000000000000000010110101011110; // input=2.779296875, output=0.35442191493
			11'd712: out = 32'b00000000000000000010110011100110; // input=2.783203125, output=0.350766542017
			11'd713: out = 32'b00000000000000000010110001101110; // input=2.787109375, output=0.347105816838
			11'd714: out = 32'b00000000000000000010101111110110; // input=2.791015625, output=0.343439795251
			11'd715: out = 32'b00000000000000000010101101111110; // input=2.794921875, output=0.339768533196
			11'd716: out = 32'b00000000000000000010101100000101; // input=2.798828125, output=0.336092086691
			11'd717: out = 32'b00000000000000000010101010001100; // input=2.802734375, output=0.332410511834
			11'd718: out = 32'b00000000000000000010101000010100; // input=2.806640625, output=0.328723864801
			11'd719: out = 32'b00000000000000000010100110011011; // input=2.810546875, output=0.325032201847
			11'd720: out = 32'b00000000000000000010100100100010; // input=2.814453125, output=0.321335579302
			11'd721: out = 32'b00000000000000000010100010101000; // input=2.818359375, output=0.31763405357
			11'd722: out = 32'b00000000000000000010100000101111; // input=2.822265625, output=0.313927681134
			11'd723: out = 32'b00000000000000000010011110110101; // input=2.826171875, output=0.310216518548
			11'd724: out = 32'b00000000000000000010011100111011; // input=2.830078125, output=0.306500622439
			11'd725: out = 32'b00000000000000000010011011000001; // input=2.833984375, output=0.302780049508
			11'd726: out = 32'b00000000000000000010011001000111; // input=2.837890625, output=0.299054856526
			11'd727: out = 32'b00000000000000000010010111001101; // input=2.841796875, output=0.295325100335
			11'd728: out = 32'b00000000000000000010010101010011; // input=2.845703125, output=0.291590837846
			11'd729: out = 32'b00000000000000000010010011011000; // input=2.849609375, output=0.28785212604
			11'd730: out = 32'b00000000000000000010010001011110; // input=2.853515625, output=0.284109021964
			11'd731: out = 32'b00000000000000000010001111100011; // input=2.857421875, output=0.280361582734
			11'd732: out = 32'b00000000000000000010001101101000; // input=2.861328125, output=0.276609865532
			11'd733: out = 32'b00000000000000000010001011101101; // input=2.865234375, output=0.272853927603
			11'd734: out = 32'b00000000000000000010001001110010; // input=2.869140625, output=0.269093826259
			11'd735: out = 32'b00000000000000000010000111110110; // input=2.873046875, output=0.265329618874
			11'd736: out = 32'b00000000000000000010000101111011; // input=2.876953125, output=0.261561362886
			11'd737: out = 32'b00000000000000000010000011111111; // input=2.880859375, output=0.257789115793
			11'd738: out = 32'b00000000000000000010000010000011; // input=2.884765625, output=0.254012935156
			11'd739: out = 32'b00000000000000000010000000001000; // input=2.888671875, output=0.250232878593
			11'd740: out = 32'b00000000000000000001111110001100; // input=2.892578125, output=0.246449003785
			11'd741: out = 32'b00000000000000000001111100010000; // input=2.896484375, output=0.242661368468
			11'd742: out = 32'b00000000000000000001111010010011; // input=2.900390625, output=0.238870030437
			11'd743: out = 32'b00000000000000000001111000010111; // input=2.904296875, output=0.235075047543
			11'd744: out = 32'b00000000000000000001110110011010; // input=2.908203125, output=0.231276477694
			11'd745: out = 32'b00000000000000000001110100011110; // input=2.912109375, output=0.22747437885
			11'd746: out = 32'b00000000000000000001110010100001; // input=2.916015625, output=0.223668809027
			11'd747: out = 32'b00000000000000000001110000100100; // input=2.919921875, output=0.219859826292
			11'd748: out = 32'b00000000000000000001101110100111; // input=2.923828125, output=0.216047488768
			11'd749: out = 32'b00000000000000000001101100101010; // input=2.927734375, output=0.212231854624
			11'd750: out = 32'b00000000000000000001101010101101; // input=2.931640625, output=0.208412982084
			11'd751: out = 32'b00000000000000000001101000110000; // input=2.935546875, output=0.204590929418
			11'd752: out = 32'b00000000000000000001100110110011; // input=2.939453125, output=0.200765754946
			11'd753: out = 32'b00000000000000000001100100110101; // input=2.943359375, output=0.196937517036
			11'd754: out = 32'b00000000000000000001100010111000; // input=2.947265625, output=0.193106274101
			11'd755: out = 32'b00000000000000000001100000111010; // input=2.951171875, output=0.189272084602
			11'd756: out = 32'b00000000000000000001011110111100; // input=2.955078125, output=0.185435007044
			11'd757: out = 32'b00000000000000000001011100111111; // input=2.958984375, output=0.181595099977
			11'd758: out = 32'b00000000000000000001011011000001; // input=2.962890625, output=0.177752421991
			11'd759: out = 32'b00000000000000000001011001000011; // input=2.966796875, output=0.173907031722
			11'd760: out = 32'b00000000000000000001010111000100; // input=2.970703125, output=0.170058987846
			11'd761: out = 32'b00000000000000000001010101000110; // input=2.974609375, output=0.166208349078
			11'd762: out = 32'b00000000000000000001010011001000; // input=2.978515625, output=0.162355174176
			11'd763: out = 32'b00000000000000000001010001001010; // input=2.982421875, output=0.158499521934
			11'd764: out = 32'b00000000000000000001001111001011; // input=2.986328125, output=0.154641451184
			11'd765: out = 32'b00000000000000000001001101001101; // input=2.990234375, output=0.150781020795
			11'd766: out = 32'b00000000000000000001001011001110; // input=2.994140625, output=0.146918289674
			11'd767: out = 32'b00000000000000000001001001010000; // input=2.998046875, output=0.14305331676
			11'd768: out = 32'b00000000000000000001000111010001; // input=3.001953125, output=0.139186161029
			11'd769: out = 32'b00000000000000000001000101010010; // input=3.005859375, output=0.135316881489
			11'd770: out = 32'b00000000000000000001000011010011; // input=3.009765625, output=0.131445537179
			11'd771: out = 32'b00000000000000000001000001010100; // input=3.013671875, output=0.127572187172
			11'd772: out = 32'b00000000000000000000111111010101; // input=3.017578125, output=0.12369689057
			11'd773: out = 32'b00000000000000000000111101010110; // input=3.021484375, output=0.119819706506
			11'd774: out = 32'b00000000000000000000111011010111; // input=3.025390625, output=0.115940694141
			11'd775: out = 32'b00000000000000000000111001011000; // input=3.029296875, output=0.112059912663
			11'd776: out = 32'b00000000000000000000110111011001; // input=3.033203125, output=0.108177421289
			11'd777: out = 32'b00000000000000000000110101011001; // input=3.037109375, output=0.10429327926
			11'd778: out = 32'b00000000000000000000110011011010; // input=3.041015625, output=0.100407545845
			11'd779: out = 32'b00000000000000000000110001011011; // input=3.044921875, output=0.0965202803338
			11'd780: out = 32'b00000000000000000000101111011011; // input=3.048828125, output=0.0926315420419
			11'd781: out = 32'b00000000000000000000101101011100; // input=3.052734375, output=0.0887413903066
			11'd782: out = 32'b00000000000000000000101011011100; // input=3.056640625, output=0.0848498844869
			11'd783: out = 32'b00000000000000000000101001011101; // input=3.060546875, output=0.0809570839624
			11'd784: out = 32'b00000000000000000000100111011101; // input=3.064453125, output=0.0770630481324
			11'd785: out = 32'b00000000000000000000100101011110; // input=3.068359375, output=0.0731678364151
			11'd786: out = 32'b00000000000000000000100011011110; // input=3.072265625, output=0.0692715082466
			11'd787: out = 32'b00000000000000000000100001011110; // input=3.076171875, output=0.0653741230801
			11'd788: out = 32'b00000000000000000000011111011110; // input=3.080078125, output=0.061475740385
			11'd789: out = 32'b00000000000000000000011101011111; // input=3.083984375, output=0.0575764196456
			11'd790: out = 32'b00000000000000000000011011011111; // input=3.087890625, output=0.053676220361
			11'd791: out = 32'b00000000000000000000011001011111; // input=3.091796875, output=0.0497752020432
			11'd792: out = 32'b00000000000000000000010111011111; // input=3.095703125, output=0.0458734242172
			11'd793: out = 32'b00000000000000000000010101011111; // input=3.099609375, output=0.0419709464191
			11'd794: out = 32'b00000000000000000000010011011111; // input=3.103515625, output=0.038067828196
			11'd795: out = 32'b00000000000000000000010001011111; // input=3.107421875, output=0.0341641291047
			11'd796: out = 32'b00000000000000000000001111100000; // input=3.111328125, output=0.0302599087108
			11'd797: out = 32'b00000000000000000000001101100000; // input=3.115234375, output=0.0263552265879
			11'd798: out = 32'b00000000000000000000001011100000; // input=3.119140625, output=0.0224501423167
			11'd799: out = 32'b00000000000000000000001001100000; // input=3.123046875, output=0.018544715484
			11'd800: out = 32'b00000000000000000000000111100000; // input=3.126953125, output=0.0146390056817
			11'd801: out = 32'b00000000000000000000000101100000; // input=3.130859375, output=0.0107330725062
			11'd802: out = 32'b00000000000000000000000011100000; // input=3.134765625, output=0.0068269755572
			11'd803: out = 32'b00000000000000000000000001100000; // input=3.138671875, output=0.00292077443696
			11'd804: out = 32'b10000000000000000000000000100000; // input=3.142578125, output=-0.000985471250699
			11'd805: out = 32'b10000000000000000000000010100000; // input=3.146484375, output=-0.00489170190128
			11'd806: out = 32'b10000000000000000000000100100000; // input=3.150390625, output=-0.00879785791051
			11'd807: out = 32'b10000000000000000000000110100000; // input=3.154296875, output=-0.0127038796752
			11'd808: out = 32'b10000000000000000000001000100000; // input=3.158203125, output=-0.0166097075944
			11'd809: out = 32'b10000000000000000000001010100000; // input=3.162109375, output=-0.0205152820699
			11'd810: out = 32'b10000000000000000000001100100000; // input=3.166015625, output=-0.0244205435074
			11'd811: out = 32'b10000000000000000000001110100000; // input=3.169921875, output=-0.0283254323174
			11'd812: out = 32'b10000000000000000000010000100000; // input=3.173828125, output=-0.0322298889162
			11'd813: out = 32'b10000000000000000000010010100000; // input=3.177734375, output=-0.0361338537266
			11'd814: out = 32'b10000000000000000000010100100000; // input=3.181640625, output=-0.0400372671788
			11'd815: out = 32'b10000000000000000000010110100000; // input=3.185546875, output=-0.0439400697116
			11'd816: out = 32'b10000000000000000000011000100000; // input=3.189453125, output=-0.0478422017729
			11'd817: out = 32'b10000000000000000000011010100000; // input=3.193359375, output=-0.0517436038212
			11'd818: out = 32'b10000000000000000000011100011111; // input=3.197265625, output=-0.0556442163256
			11'd819: out = 32'b10000000000000000000011110011111; // input=3.201171875, output=-0.0595439797679
			11'd820: out = 32'b10000000000000000000100000011111; // input=3.205078125, output=-0.0634428346422
			11'd821: out = 32'b10000000000000000000100010011111; // input=3.208984375, output=-0.0673407214569
			11'd822: out = 32'b10000000000000000000100100011110; // input=3.212890625, output=-0.0712375807351
			11'd823: out = 32'b10000000000000000000100110011110; // input=3.216796875, output=-0.0751333530155
			11'd824: out = 32'b10000000000000000000101000011110; // input=3.220703125, output=-0.0790279788533
			11'd825: out = 32'b10000000000000000000101010011101; // input=3.224609375, output=-0.0829213988214
			11'd826: out = 32'b10000000000000000000101100011101; // input=3.228515625, output=-0.086813553511
			11'd827: out = 32'b10000000000000000000101110011100; // input=3.232421875, output=-0.0907043835325
			11'd828: out = 32'b10000000000000000000110000011100; // input=3.236328125, output=-0.0945938295168
			11'd829: out = 32'b10000000000000000000110010011011; // input=3.240234375, output=-0.0984818321156
			11'd830: out = 32'b10000000000000000000110100011010; // input=3.244140625, output=-0.102368332003
			11'd831: out = 32'b10000000000000000000110110011010; // input=3.248046875, output=-0.106253269875
			11'd832: out = 32'b10000000000000000000111000011001; // input=3.251953125, output=-0.110136586453
			11'd833: out = 32'b10000000000000000000111010011000; // input=3.255859375, output=-0.114018222483
			11'd834: out = 32'b10000000000000000000111100010111; // input=3.259765625, output=-0.117898118735
			11'd835: out = 32'b10000000000000000000111110010110; // input=3.263671875, output=-0.121776216006
			11'd836: out = 32'b10000000000000000001000000010101; // input=3.267578125, output=-0.125652455122
			11'd837: out = 32'b10000000000000000001000010010100; // input=3.271484375, output=-0.129526776936
			11'd838: out = 32'b10000000000000000001000100010011; // input=3.275390625, output=-0.133399122331
			11'd839: out = 32'b10000000000000000001000110010010; // input=3.279296875, output=-0.13726943222
			11'd840: out = 32'b10000000000000000001001000010001; // input=3.283203125, output=-0.141137647546
			11'd841: out = 32'b10000000000000000001001010001111; // input=3.287109375, output=-0.145003709285
			11'd842: out = 32'b10000000000000000001001100001110; // input=3.291015625, output=-0.148867558446
			11'd843: out = 32'b10000000000000000001001110001101; // input=3.294921875, output=-0.152729136071
			11'd844: out = 32'b10000000000000000001010000001011; // input=3.298828125, output=-0.156588383237
			11'd845: out = 32'b10000000000000000001010010001001; // input=3.302734375, output=-0.160445241058
			11'd846: out = 32'b10000000000000000001010100001000; // input=3.306640625, output=-0.164299650681
			11'd847: out = 32'b10000000000000000001010110000110; // input=3.310546875, output=-0.168151553294
			11'd848: out = 32'b10000000000000000001011000000100; // input=3.314453125, output=-0.172000890121
			11'd849: out = 32'b10000000000000000001011010000010; // input=3.318359375, output=-0.175847602426
			11'd850: out = 32'b10000000000000000001011100000000; // input=3.322265625, output=-0.179691631513
			11'd851: out = 32'b10000000000000000001011101111110; // input=3.326171875, output=-0.183532918727
			11'd852: out = 32'b10000000000000000001011111111100; // input=3.330078125, output=-0.187371405454
			11'd853: out = 32'b10000000000000000001100001111001; // input=3.333984375, output=-0.191207033124
			11'd854: out = 32'b10000000000000000001100011110111; // input=3.337890625, output=-0.19503974321
			11'd855: out = 32'b10000000000000000001100101110101; // input=3.341796875, output=-0.198869477229
			11'd856: out = 32'b10000000000000000001100111110010; // input=3.345703125, output=-0.202696176745
			11'd857: out = 32'b10000000000000000001101001101111; // input=3.349609375, output=-0.206519783367
			11'd858: out = 32'b10000000000000000001101011101100; // input=3.353515625, output=-0.210340238751
			11'd859: out = 32'b10000000000000000001101101101010; // input=3.357421875, output=-0.214157484602
			11'd860: out = 32'b10000000000000000001101111100110; // input=3.361328125, output=-0.217971462672
			11'd861: out = 32'b10000000000000000001110001100011; // input=3.365234375, output=-0.221782114767
			11'd862: out = 32'b10000000000000000001110011100000; // input=3.369140625, output=-0.225589382739
			11'd863: out = 32'b10000000000000000001110101011101; // input=3.373046875, output=-0.229393208495
			11'd864: out = 32'b10000000000000000001110111011001; // input=3.376953125, output=-0.233193533993
			11'd865: out = 32'b10000000000000000001111001010110; // input=3.380859375, output=-0.236990301245
			11'd866: out = 32'b10000000000000000001111011010010; // input=3.384765625, output=-0.240783452315
			11'd867: out = 32'b10000000000000000001111101001110; // input=3.388671875, output=-0.244572929327
			11'd868: out = 32'b10000000000000000001111111001010; // input=3.392578125, output=-0.248358674457
			11'd869: out = 32'b10000000000000000010000001000110; // input=3.396484375, output=-0.252140629939
			11'd870: out = 32'b10000000000000000010000011000010; // input=3.400390625, output=-0.255918738065
			11'd871: out = 32'b10000000000000000010000100111110; // input=3.404296875, output=-0.259692941186
			11'd872: out = 32'b10000000000000000010000110111001; // input=3.408203125, output=-0.263463181712
			11'd873: out = 32'b10000000000000000010001000110101; // input=3.412109375, output=-0.267229402115
			11'd874: out = 32'b10000000000000000010001010110000; // input=3.416015625, output=-0.270991544925
			11'd875: out = 32'b10000000000000000010001100101011; // input=3.419921875, output=-0.274749552738
			11'd876: out = 32'b10000000000000000010001110100110; // input=3.423828125, output=-0.27850336821
			11'd877: out = 32'b10000000000000000010010000100001; // input=3.427734375, output=-0.282252934064
			11'd878: out = 32'b10000000000000000010010010011100; // input=3.431640625, output=-0.285998193086
			11'd879: out = 32'b10000000000000000010010100010110; // input=3.435546875, output=-0.289739088127
			11'd880: out = 32'b10000000000000000010010110010001; // input=3.439453125, output=-0.293475562106
			11'd881: out = 32'b10000000000000000010011000001011; // input=3.443359375, output=-0.297207558008
			11'd882: out = 32'b10000000000000000010011010000101; // input=3.447265625, output=-0.30093501889
			11'd883: out = 32'b10000000000000000010011011111111; // input=3.451171875, output=-0.304657887873
			11'd884: out = 32'b10000000000000000010011101111001; // input=3.455078125, output=-0.308376108151
			11'd885: out = 32'b10000000000000000010011111110011; // input=3.458984375, output=-0.31208962299
			11'd886: out = 32'b10000000000000000010100001101100; // input=3.462890625, output=-0.315798375725
			11'd887: out = 32'b10000000000000000010100011100101; // input=3.466796875, output=-0.319502309765
			11'd888: out = 32'b10000000000000000010100101011111; // input=3.470703125, output=-0.323201368593
			11'd889: out = 32'b10000000000000000010100111011000; // input=3.474609375, output=-0.326895495766
			11'd890: out = 32'b10000000000000000010101001010001; // input=3.478515625, output=-0.330584634915
			11'd891: out = 32'b10000000000000000010101011001001; // input=3.482421875, output=-0.33426872975
			11'd892: out = 32'b10000000000000000010101101000010; // input=3.486328125, output=-0.337947724056
			11'd893: out = 32'b10000000000000000010101110111010; // input=3.490234375, output=-0.341621561694
			11'd894: out = 32'b10000000000000000010110000110010; // input=3.494140625, output=-0.345290186609
			11'd895: out = 32'b10000000000000000010110010101011; // input=3.498046875, output=-0.348953542819
			11'd896: out = 32'b10000000000000000010110100100010; // input=3.501953125, output=-0.352611574428
			11'd897: out = 32'b10000000000000000010110110011010; // input=3.505859375, output=-0.356264225619
			11'd898: out = 32'b10000000000000000010111000010010; // input=3.509765625, output=-0.359911440655
			11'd899: out = 32'b10000000000000000010111010001001; // input=3.513671875, output=-0.363553163886
			11'd900: out = 32'b10000000000000000010111100000000; // input=3.517578125, output=-0.367189339743
			11'd901: out = 32'b10000000000000000010111101110111; // input=3.521484375, output=-0.370819912742
			11'd902: out = 32'b10000000000000000010111111101110; // input=3.525390625, output=-0.374444827485
			11'd903: out = 32'b10000000000000000011000001100100; // input=3.529296875, output=-0.378064028661
			11'd904: out = 32'b10000000000000000011000011011011; // input=3.533203125, output=-0.381677461046
			11'd905: out = 32'b10000000000000000011000101010001; // input=3.537109375, output=-0.385285069501
			11'd906: out = 32'b10000000000000000011000111000111; // input=3.541015625, output=-0.388886798981
			11'd907: out = 32'b10000000000000000011001000111101; // input=3.544921875, output=-0.392482594526
			11'd908: out = 32'b10000000000000000011001010110011; // input=3.548828125, output=-0.39607240127
			11'd909: out = 32'b10000000000000000011001100101000; // input=3.552734375, output=-0.399656164437
			11'd910: out = 32'b10000000000000000011001110011101; // input=3.556640625, output=-0.403233829342
			11'd911: out = 32'b10000000000000000011010000010010; // input=3.560546875, output=-0.406805341395
			11'd912: out = 32'b10000000000000000011010010000111; // input=3.564453125, output=-0.410370646099
			11'd913: out = 32'b10000000000000000011010011111100; // input=3.568359375, output=-0.413929689052
			11'd914: out = 32'b10000000000000000011010101110000; // input=3.572265625, output=-0.417482415947
			11'd915: out = 32'b10000000000000000011010111100100; // input=3.576171875, output=-0.421028772574
			11'd916: out = 32'b10000000000000000011011001011000; // input=3.580078125, output=-0.42456870482
			11'd917: out = 32'b10000000000000000011011011001100; // input=3.583984375, output=-0.42810215867
			11'd918: out = 32'b10000000000000000011011101000000; // input=3.587890625, output=-0.431629080208
			11'd919: out = 32'b10000000000000000011011110110011; // input=3.591796875, output=-0.435149415617
			11'd920: out = 32'b10000000000000000011100000100110; // input=3.595703125, output=-0.438663111181
			11'd921: out = 32'b10000000000000000011100010011001; // input=3.599609375, output=-0.442170113286
			11'd922: out = 32'b10000000000000000011100100001100; // input=3.603515625, output=-0.445670368419
			11'd923: out = 32'b10000000000000000011100101111110; // input=3.607421875, output=-0.44916382317
			11'd924: out = 32'b10000000000000000011100111110000; // input=3.611328125, output=-0.452650424234
			11'd925: out = 32'b10000000000000000011101001100010; // input=3.615234375, output=-0.45613011841
			11'd926: out = 32'b10000000000000000011101011010100; // input=3.619140625, output=-0.459602852601
			11'd927: out = 32'b10000000000000000011101101000110; // input=3.623046875, output=-0.463068573818
			11'd928: out = 32'b10000000000000000011101110110111; // input=3.626953125, output=-0.466527229179
			11'd929: out = 32'b10000000000000000011110000101000; // input=3.630859375, output=-0.469978765908
			11'd930: out = 32'b10000000000000000011110010011001; // input=3.634765625, output=-0.473423131339
			11'd931: out = 32'b10000000000000000011110100001010; // input=3.638671875, output=-0.476860272915
			11'd932: out = 32'b10000000000000000011110101111010; // input=3.642578125, output=-0.480290138191
			11'd933: out = 32'b10000000000000000011110111101010; // input=3.646484375, output=-0.48371267483
			11'd934: out = 32'b10000000000000000011111001011010; // input=3.650390625, output=-0.487127830609
			11'd935: out = 32'b10000000000000000011111011001010; // input=3.654296875, output=-0.490535553416
			11'd936: out = 32'b10000000000000000011111100111001; // input=3.658203125, output=-0.493935791254
			11'd937: out = 32'b10000000000000000011111110101000; // input=3.662109375, output=-0.49732849224
			11'd938: out = 32'b10000000000000000100000000010111; // input=3.666015625, output=-0.500713604605
			11'd939: out = 32'b10000000000000000100000010000110; // input=3.669921875, output=-0.504091076697
			11'd940: out = 32'b10000000000000000100000011110100; // input=3.673828125, output=-0.507460856978
			11'd941: out = 32'b10000000000000000100000101100011; // input=3.677734375, output=-0.510822894032
			11'd942: out = 32'b10000000000000000100000111010001; // input=3.681640625, output=-0.514177136557
			11'd943: out = 32'b10000000000000000100001000111110; // input=3.685546875, output=-0.517523533371
			11'd944: out = 32'b10000000000000000100001010101100; // input=3.689453125, output=-0.520862033412
			11'd945: out = 32'b10000000000000000100001100011001; // input=3.693359375, output=-0.52419258574
			11'd946: out = 32'b10000000000000000100001110000110; // input=3.697265625, output=-0.527515139534
			11'd947: out = 32'b10000000000000000100001111110010; // input=3.701171875, output=-0.530829644096
			11'd948: out = 32'b10000000000000000100010001011111; // input=3.705078125, output=-0.534136048851
			11'd949: out = 32'b10000000000000000100010011001011; // input=3.708984375, output=-0.537434303347
			11'd950: out = 32'b10000000000000000100010100110110; // input=3.712890625, output=-0.540724357256
			11'd951: out = 32'b10000000000000000100010110100010; // input=3.716796875, output=-0.544006160377
			11'd952: out = 32'b10000000000000000100011000001101; // input=3.720703125, output=-0.547279662634
			11'd953: out = 32'b10000000000000000100011001111000; // input=3.724609375, output=-0.550544814076
			11'd954: out = 32'b10000000000000000100011011100011; // input=3.728515625, output=-0.553801564881
			11'd955: out = 32'b10000000000000000100011101001101; // input=3.732421875, output=-0.557049865356
			11'd956: out = 32'b10000000000000000100011110111000; // input=3.736328125, output=-0.560289665936
			11'd957: out = 32'b10000000000000000100100000100001; // input=3.740234375, output=-0.563520917184
			11'd958: out = 32'b10000000000000000100100010001011; // input=3.744140625, output=-0.566743569797
			11'd959: out = 32'b10000000000000000100100011110100; // input=3.748046875, output=-0.5699575746
			11'd960: out = 32'b10000000000000000100100101011101; // input=3.751953125, output=-0.573162882552
			11'd961: out = 32'b10000000000000000100100111000110; // input=3.755859375, output=-0.576359444743
			11'd962: out = 32'b10000000000000000100101000101111; // input=3.759765625, output=-0.579547212398
			11'd963: out = 32'b10000000000000000100101010010111; // input=3.763671875, output=-0.582726136876
			11'd964: out = 32'b10000000000000000100101011111111; // input=3.767578125, output=-0.58589616967
			11'd965: out = 32'b10000000000000000100101101100110; // input=3.771484375, output=-0.58905726241
			11'd966: out = 32'b10000000000000000100101111001110; // input=3.775390625, output=-0.59220936686
			11'd967: out = 32'b10000000000000000100110000110101; // input=3.779296875, output=-0.595352434924
			11'd968: out = 32'b10000000000000000100110010011011; // input=3.783203125, output=-0.598486418642
			11'd969: out = 32'b10000000000000000100110100000010; // input=3.787109375, output=-0.601611270194
			11'd970: out = 32'b10000000000000000100110101101000; // input=3.791015625, output=-0.604726941898
			11'd971: out = 32'b10000000000000000100110111001101; // input=3.794921875, output=-0.607833386213
			11'd972: out = 32'b10000000000000000100111000110011; // input=3.798828125, output=-0.610930555738
			11'd973: out = 32'b10000000000000000100111010011000; // input=3.802734375, output=-0.614018403215
			11'd974: out = 32'b10000000000000000100111011111101; // input=3.806640625, output=-0.617096881526
			11'd975: out = 32'b10000000000000000100111101100010; // input=3.810546875, output=-0.620165943698
			11'd976: out = 32'b10000000000000000100111111000110; // input=3.814453125, output=-0.623225542901
			11'd977: out = 32'b10000000000000000101000000101010; // input=3.818359375, output=-0.626275632449
			11'd978: out = 32'b10000000000000000101000010001101; // input=3.822265625, output=-0.629316165801
			11'd979: out = 32'b10000000000000000101000011110001; // input=3.826171875, output=-0.632347096563
			11'd980: out = 32'b10000000000000000101000101010100; // input=3.830078125, output=-0.635368378486
			11'd981: out = 32'b10000000000000000101000110110110; // input=3.833984375, output=-0.638379965469
			11'd982: out = 32'b10000000000000000101001000011001; // input=3.837890625, output=-0.64138181156
			11'd983: out = 32'b10000000000000000101001001111011; // input=3.841796875, output=-0.644373870953
			11'd984: out = 32'b10000000000000000101001011011101; // input=3.845703125, output=-0.647356097993
			11'd985: out = 32'b10000000000000000101001100111110; // input=3.849609375, output=-0.650328447176
			11'd986: out = 32'b10000000000000000101001110011111; // input=3.853515625, output=-0.653290873148
			11'd987: out = 32'b10000000000000000101010000000000; // input=3.857421875, output=-0.656243330704
			11'd988: out = 32'b10000000000000000101010001100000; // input=3.861328125, output=-0.659185774794
			11'd989: out = 32'b10000000000000000101010011000000; // input=3.865234375, output=-0.662118160521
			11'd990: out = 32'b10000000000000000101010100100000; // input=3.869140625, output=-0.665040443139
			11'd991: out = 32'b10000000000000000101010101111111; // input=3.873046875, output=-0.667952578058
			11'd992: out = 32'b10000000000000000101010111011111; // input=3.876953125, output=-0.670854520842
			11'd993: out = 32'b10000000000000000101011000111101; // input=3.880859375, output=-0.673746227212
			11'd994: out = 32'b10000000000000000101011010011100; // input=3.884765625, output=-0.676627653043
			11'd995: out = 32'b10000000000000000101011011111010; // input=3.888671875, output=-0.679498754369
			11'd996: out = 32'b10000000000000000101011101011000; // input=3.892578125, output=-0.68235948738
			11'd997: out = 32'b10000000000000000101011110110101; // input=3.896484375, output=-0.685209808425
			11'd998: out = 32'b10000000000000000101100000010010; // input=3.900390625, output=-0.688049674011
			11'd999: out = 32'b10000000000000000101100001101111; // input=3.904296875, output=-0.690879040805
			11'd1000: out = 32'b10000000000000000101100011001011; // input=3.908203125, output=-0.693697865636
			11'd1001: out = 32'b10000000000000000101100100100111; // input=3.912109375, output=-0.69650610549
			11'd1002: out = 32'b10000000000000000101100110000011; // input=3.916015625, output=-0.699303717518
			11'd1003: out = 32'b10000000000000000101100111011110; // input=3.919921875, output=-0.702090659032
			11'd1004: out = 32'b10000000000000000101101000111001; // input=3.923828125, output=-0.704866887506
			11'd1005: out = 32'b10000000000000000101101010010100; // input=3.927734375, output=-0.707632360579
			11'd1006: out = 32'b10000000000000000101101011101110; // input=3.931640625, output=-0.710387036053
			11'd1007: out = 32'b10000000000000000101101101001000; // input=3.935546875, output=-0.713130871894
			11'd1008: out = 32'b10000000000000000101101110100001; // input=3.939453125, output=-0.715863826236
			11'd1009: out = 32'b10000000000000000101101111111011; // input=3.943359375, output=-0.718585857376
			11'd1010: out = 32'b10000000000000000101110001010011; // input=3.947265625, output=-0.72129692378
			11'd1011: out = 32'b10000000000000000101110010101100; // input=3.951171875, output=-0.723996984081
			11'd1012: out = 32'b10000000000000000101110100000100; // input=3.955078125, output=-0.726685997079
			11'd1013: out = 32'b10000000000000000101110101011100; // input=3.958984375, output=-0.729363921742
			11'd1014: out = 32'b10000000000000000101110110110011; // input=3.962890625, output=-0.732030717209
			11'd1015: out = 32'b10000000000000000101111000001010; // input=3.966796875, output=-0.734686342788
			11'd1016: out = 32'b10000000000000000101111001100001; // input=3.970703125, output=-0.737330757958
			11'd1017: out = 32'b10000000000000000101111010110111; // input=3.974609375, output=-0.739963922367
			11'd1018: out = 32'b10000000000000000101111100001101; // input=3.978515625, output=-0.742585795837
			11'd1019: out = 32'b10000000000000000101111101100011; // input=3.982421875, output=-0.745196338362
			11'd1020: out = 32'b10000000000000000101111110111000; // input=3.986328125, output=-0.747795510107
			11'd1021: out = 32'b10000000000000000110000000001101; // input=3.990234375, output=-0.750383271413
			11'd1022: out = 32'b10000000000000000110000001100001; // input=3.994140625, output=-0.752959582793
			11'd1023: out = 32'b10000000000000000110000010110101; // input=3.998046875, output=-0.755524404937
			11'd1024: out = 32'b10000000000000000000000001000000; // input=-0.001953125, output=-0.00195312375824
			11'd1025: out = 32'b10000000000000000000000011000000; // input=-0.005859375, output=-0.00585934147244
			11'd1026: out = 32'b10000000000000000000000101000000; // input=-0.009765625, output=-0.00976546978031
			11'd1027: out = 32'b10000000000000000000000111000000; // input=-0.013671875, output=-0.0136714490791
			11'd1028: out = 32'b10000000000000000000001001000000; // input=-0.017578125, output=-0.0175772197684
			11'd1029: out = 32'b10000000000000000000001011000000; // input=-0.021484375, output=-0.021482722251
			11'd1030: out = 32'b10000000000000000000001101000000; // input=-0.025390625, output=-0.0253878969337
			11'd1031: out = 32'b10000000000000000000001111000000; // input=-0.029296875, output=-0.0292926842283
			11'd1032: out = 32'b10000000000000000000010001000000; // input=-0.033203125, output=-0.0331970245525
			11'd1033: out = 32'b10000000000000000000010011000000; // input=-0.037109375, output=-0.0371008583311
			11'd1034: out = 32'b10000000000000000000010101000000; // input=-0.041015625, output=-0.0410041259961
			11'd1035: out = 32'b10000000000000000000010111000000; // input=-0.044921875, output=-0.0449067679887
			11'd1036: out = 32'b10000000000000000000011000111111; // input=-0.048828125, output=-0.0488087247592
			11'd1037: out = 32'b10000000000000000000011010111111; // input=-0.052734375, output=-0.0527099367686
			11'd1038: out = 32'b10000000000000000000011100111111; // input=-0.056640625, output=-0.0566103444893
			11'd1039: out = 32'b10000000000000000000011110111111; // input=-0.060546875, output=-0.0605098884057
			11'd1040: out = 32'b10000000000000000000100000111111; // input=-0.064453125, output=-0.0644085090157
			11'd1041: out = 32'b10000000000000000000100010111110; // input=-0.068359375, output=-0.0683061468311
			11'd1042: out = 32'b10000000000000000000100100111110; // input=-0.072265625, output=-0.0722027423787
			11'd1043: out = 32'b10000000000000000000100110111110; // input=-0.076171875, output=-0.0760982362014
			11'd1044: out = 32'b10000000000000000000101000111101; // input=-0.080078125, output=-0.0799925688585
			11'd1045: out = 32'b10000000000000000000101010111101; // input=-0.083984375, output=-0.0838856809275
			11'd1046: out = 32'b10000000000000000000101100111100; // input=-0.087890625, output=-0.0877775130042
			11'd1047: out = 32'b10000000000000000000101110111100; // input=-0.091796875, output=-0.091668005704
			11'd1048: out = 32'b10000000000000000000110000111011; // input=-0.095703125, output=-0.0955570996629
			11'd1049: out = 32'b10000000000000000000110010111011; // input=-0.099609375, output=-0.099444735538
			11'd1050: out = 32'b10000000000000000000110100111010; // input=-0.103515625, output=-0.103330854009
			11'd1051: out = 32'b10000000000000000000110110111001; // input=-0.107421875, output=-0.107215395778
			11'd1052: out = 32'b10000000000000000000111000111000; // input=-0.111328125, output=-0.111098301572
			11'd1053: out = 32'b10000000000000000000111010111000; // input=-0.115234375, output=-0.114979512142
			11'd1054: out = 32'b10000000000000000000111100110111; // input=-0.119140625, output=-0.118858968267
			11'd1055: out = 32'b10000000000000000000111110110110; // input=-0.123046875, output=-0.12273661075
			11'd1056: out = 32'b10000000000000000001000000110101; // input=-0.126953125, output=-0.126612380424
			11'd1057: out = 32'b10000000000000000001000010110100; // input=-0.130859375, output=-0.130486218148
			11'd1058: out = 32'b10000000000000000001000100110011; // input=-0.134765625, output=-0.134358064813
			11'd1059: out = 32'b10000000000000000001000110110001; // input=-0.138671875, output=-0.13822786134
			11'd1060: out = 32'b10000000000000000001001000110000; // input=-0.142578125, output=-0.142095548679
			11'd1061: out = 32'b10000000000000000001001010101111; // input=-0.146484375, output=-0.145961067815
			11'd1062: out = 32'b10000000000000000001001100101101; // input=-0.150390625, output=-0.149824359765
			11'd1063: out = 32'b10000000000000000001001110101100; // input=-0.154296875, output=-0.153685365579
			11'd1064: out = 32'b10000000000000000001010000101010; // input=-0.158203125, output=-0.157544026344
			11'd1065: out = 32'b10000000000000000001010010101001; // input=-0.162109375, output=-0.161400283181
			11'd1066: out = 32'b10000000000000000001010100100111; // input=-0.166015625, output=-0.165254077248
			11'd1067: out = 32'b10000000000000000001010110100101; // input=-0.169921875, output=-0.169105349741
			11'd1068: out = 32'b10000000000000000001011000100011; // input=-0.173828125, output=-0.172954041894
			11'd1069: out = 32'b10000000000000000001011010100001; // input=-0.177734375, output=-0.176800094982
			11'd1070: out = 32'b10000000000000000001011100011111; // input=-0.181640625, output=-0.180643450318
			11'd1071: out = 32'b10000000000000000001011110011101; // input=-0.185546875, output=-0.184484049257
			11'd1072: out = 32'b10000000000000000001100000011011; // input=-0.189453125, output=-0.188321833196
			11'd1073: out = 32'b10000000000000000001100010011001; // input=-0.193359375, output=-0.192156743576
			11'd1074: out = 32'b10000000000000000001100100010110; // input=-0.197265625, output=-0.19598872188
			11'd1075: out = 32'b10000000000000000001100110010100; // input=-0.201171875, output=-0.199817709638
			11'd1076: out = 32'b10000000000000000001101000010001; // input=-0.205078125, output=-0.203643648423
			11'd1077: out = 32'b10000000000000000001101010001110; // input=-0.208984375, output=-0.207466479857
			11'd1078: out = 32'b10000000000000000001101100001011; // input=-0.212890625, output=-0.211286145607
			11'd1079: out = 32'b10000000000000000001101110001000; // input=-0.216796875, output=-0.215102587391
			11'd1080: out = 32'b10000000000000000001110000000101; // input=-0.220703125, output=-0.218915746974
			11'd1081: out = 32'b10000000000000000001110010000010; // input=-0.224609375, output=-0.222725566172
			11'd1082: out = 32'b10000000000000000001110011111111; // input=-0.228515625, output=-0.226531986852
			11'd1083: out = 32'b10000000000000000001110101111100; // input=-0.232421875, output=-0.230334950932
			11'd1084: out = 32'b10000000000000000001110111111000; // input=-0.236328125, output=-0.234134400385
			11'd1085: out = 32'b10000000000000000001111001110100; // input=-0.240234375, output=-0.237930277234
			11'd1086: out = 32'b10000000000000000001111011110001; // input=-0.244140625, output=-0.241722523561
			11'd1087: out = 32'b10000000000000000001111101101101; // input=-0.248046875, output=-0.245511081499
			11'd1088: out = 32'b10000000000000000001111111101001; // input=-0.251953125, output=-0.24929589324
			11'd1089: out = 32'b10000000000000000010000001100101; // input=-0.255859375, output=-0.253076901032
			11'd1090: out = 32'b10000000000000000010000011100001; // input=-0.259765625, output=-0.256854047182
			11'd1091: out = 32'b10000000000000000010000101011100; // input=-0.263671875, output=-0.260627274056
			11'd1092: out = 32'b10000000000000000010000111011000; // input=-0.267578125, output=-0.264396524078
			11'd1093: out = 32'b10000000000000000010001001010011; // input=-0.271484375, output=-0.268161739734
			11'd1094: out = 32'b10000000000000000010001011001110; // input=-0.275390625, output=-0.271922863572
			11'd1095: out = 32'b10000000000000000010001101001001; // input=-0.279296875, output=-0.275679838202
			11'd1096: out = 32'b10000000000000000010001111000100; // input=-0.283203125, output=-0.279432606296
			11'd1097: out = 32'b10000000000000000010010000111111; // input=-0.287109375, output=-0.283181110593
			11'd1098: out = 32'b10000000000000000010010010111010; // input=-0.291015625, output=-0.286925293895
			11'd1099: out = 32'b10000000000000000010010100110101; // input=-0.294921875, output=-0.290665099069
			11'd1100: out = 32'b10000000000000000010010110101111; // input=-0.298828125, output=-0.294400469052
			11'd1101: out = 32'b10000000000000000010011000101001; // input=-0.302734375, output=-0.298131346846
			11'd1102: out = 32'b10000000000000000010011010100011; // input=-0.306640625, output=-0.301857675522
			11'd1103: out = 32'b10000000000000000010011100011101; // input=-0.310546875, output=-0.305579398221
			11'd1104: out = 32'b10000000000000000010011110010111; // input=-0.314453125, output=-0.309296458155
			11'd1105: out = 32'b10000000000000000010100000010001; // input=-0.318359375, output=-0.313008798605
			11'd1106: out = 32'b10000000000000000010100010001010; // input=-0.322265625, output=-0.316716362927
			11'd1107: out = 32'b10000000000000000010100100000011; // input=-0.326171875, output=-0.320419094546
			11'd1108: out = 32'b10000000000000000010100101111101; // input=-0.330078125, output=-0.324116936964
			11'd1109: out = 32'b10000000000000000010100111110110; // input=-0.333984375, output=-0.327809833756
			11'd1110: out = 32'b10000000000000000010101001101111; // input=-0.337890625, output=-0.331497728574
			11'd1111: out = 32'b10000000000000000010101011100111; // input=-0.341796875, output=-0.335180565144
			11'd1112: out = 32'b10000000000000000010101101100000; // input=-0.345703125, output=-0.338858287271
			11'd1113: out = 32'b10000000000000000010101111011000; // input=-0.349609375, output=-0.342530838838
			11'd1114: out = 32'b10000000000000000010110001010000; // input=-0.353515625, output=-0.346198163805
			11'd1115: out = 32'b10000000000000000010110011001000; // input=-0.357421875, output=-0.349860206215
			11'd1116: out = 32'b10000000000000000010110101000000; // input=-0.361328125, output=-0.353516910188
			11'd1117: out = 32'b10000000000000000010110110111000; // input=-0.365234375, output=-0.357168219928
			11'd1118: out = 32'b10000000000000000010111000101111; // input=-0.369140625, output=-0.36081407972
			11'd1119: out = 32'b10000000000000000010111010100110; // input=-0.373046875, output=-0.364454433933
			11'd1120: out = 32'b10000000000000000010111100011110; // input=-0.376953125, output=-0.36808922702
			11'd1121: out = 32'b10000000000000000010111110010100; // input=-0.380859375, output=-0.371718403519
			11'd1122: out = 32'b10000000000000000011000000001011; // input=-0.384765625, output=-0.375341908052
			11'd1123: out = 32'b10000000000000000011000010000010; // input=-0.388671875, output=-0.378959685329
			11'd1124: out = 32'b10000000000000000011000011111000; // input=-0.392578125, output=-0.382571680148
			11'd1125: out = 32'b10000000000000000011000101101110; // input=-0.396484375, output=-0.386177837393
			11'd1126: out = 32'b10000000000000000011000111100100; // input=-0.400390625, output=-0.38977810204
			11'd1127: out = 32'b10000000000000000011001001011010; // input=-0.404296875, output=-0.393372419153
			11'd1128: out = 32'b10000000000000000011001011010000; // input=-0.408203125, output=-0.396960733886
			11'd1129: out = 32'b10000000000000000011001101000101; // input=-0.412109375, output=-0.400542991487
			11'd1130: out = 32'b10000000000000000011001110111010; // input=-0.416015625, output=-0.404119137295
			11'd1131: out = 32'b10000000000000000011010000101111; // input=-0.419921875, output=-0.407689116742
			11'd1132: out = 32'b10000000000000000011010010100100; // input=-0.423828125, output=-0.411252875354
			11'd1133: out = 32'b10000000000000000011010100011001; // input=-0.427734375, output=-0.414810358754
			11'd1134: out = 32'b10000000000000000011010110001101; // input=-0.431640625, output=-0.418361512658
			11'd1135: out = 32'b10000000000000000011011000000001; // input=-0.435546875, output=-0.42190628288
			11'd1136: out = 32'b10000000000000000011011001110101; // input=-0.439453125, output=-0.425444615332
			11'd1137: out = 32'b10000000000000000011011011101001; // input=-0.443359375, output=-0.428976456021
			11'd1138: out = 32'b10000000000000000011011101011100; // input=-0.447265625, output=-0.432501751058
			11'd1139: out = 32'b10000000000000000011011111010000; // input=-0.451171875, output=-0.436020446651
			11'd1140: out = 32'b10000000000000000011100001000011; // input=-0.455078125, output=-0.439532489107
			11'd1141: out = 32'b10000000000000000011100010110101; // input=-0.458984375, output=-0.443037824839
			11'd1142: out = 32'b10000000000000000011100100101000; // input=-0.462890625, output=-0.446536400359
			11'd1143: out = 32'b10000000000000000011100110011011; // input=-0.466796875, output=-0.450028162283
			11'd1144: out = 32'b10000000000000000011101000001101; // input=-0.470703125, output=-0.45351305733
			11'd1145: out = 32'b10000000000000000011101001111111; // input=-0.474609375, output=-0.456991032326
			11'd1146: out = 32'b10000000000000000011101011110000; // input=-0.478515625, output=-0.460462034202
			11'd1147: out = 32'b10000000000000000011101101100010; // input=-0.482421875, output=-0.463926009993
			11'd1148: out = 32'b10000000000000000011101111010011; // input=-0.486328125, output=-0.467382906844
			11'd1149: out = 32'b10000000000000000011110001000100; // input=-0.490234375, output=-0.470832672007
			11'd1150: out = 32'b10000000000000000011110010110101; // input=-0.494140625, output=-0.474275252843
			11'd1151: out = 32'b10000000000000000011110100100110; // input=-0.498046875, output=-0.477710596821
			11'd1152: out = 32'b10000000000000000011110110010110; // input=-0.501953125, output=-0.481138651524
			11'd1153: out = 32'b10000000000000000011111000000110; // input=-0.505859375, output=-0.484559364643
			11'd1154: out = 32'b10000000000000000011111001110110; // input=-0.509765625, output=-0.487972683983
			11'd1155: out = 32'b10000000000000000011111011100101; // input=-0.513671875, output=-0.491378557459
			11'd1156: out = 32'b10000000000000000011111101010101; // input=-0.517578125, output=-0.494776933103
			11'd1157: out = 32'b10000000000000000011111111000100; // input=-0.521484375, output=-0.49816775906
			11'd1158: out = 32'b10000000000000000100000000110011; // input=-0.525390625, output=-0.50155098359
			11'd1159: out = 32'b10000000000000000100000010100001; // input=-0.529296875, output=-0.504926555069
			11'd1160: out = 32'b10000000000000000100000100010000; // input=-0.533203125, output=-0.50829442199
			11'd1161: out = 32'b10000000000000000100000101111110; // input=-0.537109375, output=-0.511654532964
			11'd1162: out = 32'b10000000000000000100000111101100; // input=-0.541015625, output=-0.515006836719
			11'd1163: out = 32'b10000000000000000100001001011001; // input=-0.544921875, output=-0.518351282103
			11'd1164: out = 32'b10000000000000000100001011000111; // input=-0.548828125, output=-0.521687818084
			11'd1165: out = 32'b10000000000000000100001100110100; // input=-0.552734375, output=-0.525016393751
			11'd1166: out = 32'b10000000000000000100001110100001; // input=-0.556640625, output=-0.528336958314
			11'd1167: out = 32'b10000000000000000100010000001101; // input=-0.560546875, output=-0.531649461105
			11'd1168: out = 32'b10000000000000000100010001111001; // input=-0.564453125, output=-0.534953851579
			11'd1169: out = 32'b10000000000000000100010011100101; // input=-0.568359375, output=-0.538250079316
			11'd1170: out = 32'b10000000000000000100010101010001; // input=-0.572265625, output=-0.541538094019
			11'd1171: out = 32'b10000000000000000100010110111101; // input=-0.576171875, output=-0.544817845516
			11'd1172: out = 32'b10000000000000000100011000101000; // input=-0.580078125, output=-0.548089283764
			11'd1173: out = 32'b10000000000000000100011010010011; // input=-0.583984375, output=-0.551352358843
			11'd1174: out = 32'b10000000000000000100011011111101; // input=-0.587890625, output=-0.554607020964
			11'd1175: out = 32'b10000000000000000100011101101000; // input=-0.591796875, output=-0.557853220464
			11'd1176: out = 32'b10000000000000000100011111010010; // input=-0.595703125, output=-0.561090907811
			11'd1177: out = 32'b10000000000000000100100000111100; // input=-0.599609375, output=-0.5643200336
			11'd1178: out = 32'b10000000000000000100100010100101; // input=-0.603515625, output=-0.56754054856
			11'd1179: out = 32'b10000000000000000100100100001110; // input=-0.607421875, output=-0.570752403549
			11'd1180: out = 32'b10000000000000000100100101110111; // input=-0.611328125, output=-0.573955549559
			11'd1181: out = 32'b10000000000000000100100111100000; // input=-0.615234375, output=-0.577149937714
			11'd1182: out = 32'b10000000000000000100101001001000; // input=-0.619140625, output=-0.58033551927
			11'd1183: out = 32'b10000000000000000100101010110001; // input=-0.623046875, output=-0.583512245621
			11'd1184: out = 32'b10000000000000000100101100011000; // input=-0.626953125, output=-0.586680068292
			11'd1185: out = 32'b10000000000000000100101110000000; // input=-0.630859375, output=-0.589838938948
			11'd1186: out = 32'b10000000000000000100101111100111; // input=-0.634765625, output=-0.592988809387
			11'd1187: out = 32'b10000000000000000100110001001110; // input=-0.638671875, output=-0.596129631546
			11'd1188: out = 32'b10000000000000000100110010110101; // input=-0.642578125, output=-0.599261357501
			11'd1189: out = 32'b10000000000000000100110100011011; // input=-0.646484375, output=-0.602383939464
			11'd1190: out = 32'b10000000000000000100110110000001; // input=-0.650390625, output=-0.60549732979
			11'd1191: out = 32'b10000000000000000100110111100111; // input=-0.654296875, output=-0.608601480971
			11'd1192: out = 32'b10000000000000000100111001001100; // input=-0.658203125, output=-0.611696345643
			11'd1193: out = 32'b10000000000000000100111010110001; // input=-0.662109375, output=-0.614781876581
			11'd1194: out = 32'b10000000000000000100111100010110; // input=-0.666015625, output=-0.617858026704
			11'd1195: out = 32'b10000000000000000100111101111010; // input=-0.669921875, output=-0.620924749074
			11'd1196: out = 32'b10000000000000000100111111011111; // input=-0.673828125, output=-0.623981996896
			11'd1197: out = 32'b10000000000000000101000001000011; // input=-0.677734375, output=-0.62702972352
			11'd1198: out = 32'b10000000000000000101000010100110; // input=-0.681640625, output=-0.630067882443
			11'd1199: out = 32'b10000000000000000101000100001001; // input=-0.685546875, output=-0.633096427304
			11'd1200: out = 32'b10000000000000000101000101101100; // input=-0.689453125, output=-0.636115311893
			11'd1201: out = 32'b10000000000000000101000111001111; // input=-0.693359375, output=-0.639124490145
			11'd1202: out = 32'b10000000000000000101001000110001; // input=-0.697265625, output=-0.642123916144
			11'd1203: out = 32'b10000000000000000101001010010011; // input=-0.701171875, output=-0.645113544122
			11'd1204: out = 32'b10000000000000000101001011110101; // input=-0.705078125, output=-0.64809332846
			11'd1205: out = 32'b10000000000000000101001101010110; // input=-0.708984375, output=-0.651063223692
			11'd1206: out = 32'b10000000000000000101001110110111; // input=-0.712890625, output=-0.6540231845
			11'd1207: out = 32'b10000000000000000101010000011000; // input=-0.716796875, output=-0.65697316572
			11'd1208: out = 32'b10000000000000000101010001111000; // input=-0.720703125, output=-0.659913122336
			11'd1209: out = 32'b10000000000000000101010011011000; // input=-0.724609375, output=-0.662843009491
			11'd1210: out = 32'b10000000000000000101010100111000; // input=-0.728515625, output=-0.665762782477
			11'd1211: out = 32'b10000000000000000101010110010111; // input=-0.732421875, output=-0.668672396741
			11'd1212: out = 32'b10000000000000000101010111110110; // input=-0.736328125, output=-0.671571807888
			11'd1213: out = 32'b10000000000000000101011001010101; // input=-0.740234375, output=-0.674460971675
			11'd1214: out = 32'b10000000000000000101011010110011; // input=-0.744140625, output=-0.677339844018
			11'd1215: out = 32'b10000000000000000101011100010001; // input=-0.748046875, output=-0.680208380988
			11'd1216: out = 32'b10000000000000000101011101101111; // input=-0.751953125, output=-0.683066538814
			11'd1217: out = 32'b10000000000000000101011111001100; // input=-0.755859375, output=-0.685914273886
			11'd1218: out = 32'b10000000000000000101100000101001; // input=-0.759765625, output=-0.68875154275
			11'd1219: out = 32'b10000000000000000101100010000110; // input=-0.763671875, output=-0.691578302113
			11'd1220: out = 32'b10000000000000000101100011100010; // input=-0.767578125, output=-0.694394508842
			11'd1221: out = 32'b10000000000000000101100100111110; // input=-0.771484375, output=-0.697200119965
			11'd1222: out = 32'b10000000000000000101100110011001; // input=-0.775390625, output=-0.699995092672
			11'd1223: out = 32'b10000000000000000101100111110101; // input=-0.779296875, output=-0.702779384315
			11'd1224: out = 32'b10000000000000000101101001010000; // input=-0.783203125, output=-0.705552952409
			11'd1225: out = 32'b10000000000000000101101010101010; // input=-0.787109375, output=-0.708315754633
			11'd1226: out = 32'b10000000000000000101101100000100; // input=-0.791015625, output=-0.711067748831
			11'd1227: out = 32'b10000000000000000101101101011110; // input=-0.794921875, output=-0.713808893009
			11'd1228: out = 32'b10000000000000000101101110111000; // input=-0.798828125, output=-0.716539145342
			11'd1229: out = 32'b10000000000000000101110000010001; // input=-0.802734375, output=-0.719258464169
			11'd1230: out = 32'b10000000000000000101110001101001; // input=-0.806640625, output=-0.721966807997
			11'd1231: out = 32'b10000000000000000101110011000010; // input=-0.810546875, output=-0.7246641355
			11'd1232: out = 32'b10000000000000000101110100011010; // input=-0.814453125, output=-0.727350405519
			11'd1233: out = 32'b10000000000000000101110101110001; // input=-0.818359375, output=-0.730025577067
			11'd1234: out = 32'b10000000000000000101110111001001; // input=-0.822265625, output=-0.732689609322
			11'd1235: out = 32'b10000000000000000101111000100000; // input=-0.826171875, output=-0.735342461635
			11'd1236: out = 32'b10000000000000000101111001110110; // input=-0.830078125, output=-0.737984093527
			11'd1237: out = 32'b10000000000000000101111011001100; // input=-0.833984375, output=-0.740614464689
			11'd1238: out = 32'b10000000000000000101111100100010; // input=-0.837890625, output=-0.743233534986
			11'd1239: out = 32'b10000000000000000101111101111000; // input=-0.841796875, output=-0.745841264454
			11'd1240: out = 32'b10000000000000000101111111001101; // input=-0.845703125, output=-0.748437613302
			11'd1241: out = 32'b10000000000000000110000000100010; // input=-0.849609375, output=-0.751022541912
			11'd1242: out = 32'b10000000000000000110000001110110; // input=-0.853515625, output=-0.753596010843
			11'd1243: out = 32'b10000000000000000110000011001010; // input=-0.857421875, output=-0.756157980826
			11'd1244: out = 32'b10000000000000000110000100011101; // input=-0.861328125, output=-0.758708412768
			11'd1245: out = 32'b10000000000000000110000101110001; // input=-0.865234375, output=-0.761247267753
			11'd1246: out = 32'b10000000000000000110000111000011; // input=-0.869140625, output=-0.763774507042
			11'd1247: out = 32'b10000000000000000110001000010110; // input=-0.873046875, output=-0.766290092071
			11'd1248: out = 32'b10000000000000000110001001101000; // input=-0.876953125, output=-0.768793984456
			11'd1249: out = 32'b10000000000000000110001010111010; // input=-0.880859375, output=-0.771286145991
			11'd1250: out = 32'b10000000000000000110001100001011; // input=-0.884765625, output=-0.773766538648
			11'd1251: out = 32'b10000000000000000110001101011100; // input=-0.888671875, output=-0.77623512458
			11'd1252: out = 32'b10000000000000000110001110101100; // input=-0.892578125, output=-0.778691866119
			11'd1253: out = 32'b10000000000000000110001111111100; // input=-0.896484375, output=-0.781136725778
			11'd1254: out = 32'b10000000000000000110010001001100; // input=-0.900390625, output=-0.783569666252
			11'd1255: out = 32'b10000000000000000110010010011011; // input=-0.904296875, output=-0.785990650417
			11'd1256: out = 32'b10000000000000000110010011101010; // input=-0.908203125, output=-0.788399641331
			11'd1257: out = 32'b10000000000000000110010100111001; // input=-0.912109375, output=-0.790796602237
			11'd1258: out = 32'b10000000000000000110010110000111; // input=-0.916015625, output=-0.79318149656
			11'd1259: out = 32'b10000000000000000110010111010101; // input=-0.919921875, output=-0.795554287909
			11'd1260: out = 32'b10000000000000000110011000100010; // input=-0.923828125, output=-0.797914940078
			11'd1261: out = 32'b10000000000000000110011001101111; // input=-0.927734375, output=-0.800263417047
			11'd1262: out = 32'b10000000000000000110011010111100; // input=-0.931640625, output=-0.802599682981
			11'd1263: out = 32'b10000000000000000110011100001000; // input=-0.935546875, output=-0.804923702231
			11'd1264: out = 32'b10000000000000000110011101010011; // input=-0.939453125, output=-0.807235439336
			11'd1265: out = 32'b10000000000000000110011110011111; // input=-0.943359375, output=-0.809534859021
			11'd1266: out = 32'b10000000000000000110011111101010; // input=-0.947265625, output=-0.8118219262
			11'd1267: out = 32'b10000000000000000110100000110100; // input=-0.951171875, output=-0.814096605976
			11'd1268: out = 32'b10000000000000000110100001111110; // input=-0.955078125, output=-0.816358863639
			11'd1269: out = 32'b10000000000000000110100011001000; // input=-0.958984375, output=-0.81860866467
			11'd1270: out = 32'b10000000000000000110100100010001; // input=-0.962890625, output=-0.82084597474
			11'd1271: out = 32'b10000000000000000110100101011010; // input=-0.966796875, output=-0.82307075971
			11'd1272: out = 32'b10000000000000000110100110100011; // input=-0.970703125, output=-0.825282985633
			11'd1273: out = 32'b10000000000000000110100111101011; // input=-0.974609375, output=-0.827482618753
			11'd1274: out = 32'b10000000000000000110101000110011; // input=-0.978515625, output=-0.829669625507
			11'd1275: out = 32'b10000000000000000110101001111010; // input=-0.982421875, output=-0.831843972523
			11'd1276: out = 32'b10000000000000000110101011000001; // input=-0.986328125, output=-0.834005626623
			11'd1277: out = 32'b10000000000000000110101100000111; // input=-0.990234375, output=-0.836154554823
			11'd1278: out = 32'b10000000000000000110101101001101; // input=-0.994140625, output=-0.838290724334
			11'd1279: out = 32'b10000000000000000110101110010011; // input=-0.998046875, output=-0.84041410256
			11'd1280: out = 32'b10000000000000000110101111011000; // input=-1.001953125, output=-0.8425246571
			11'd1281: out = 32'b10000000000000000110110000011101; // input=-1.005859375, output=-0.844622355751
			11'd1282: out = 32'b10000000000000000110110001100001; // input=-1.009765625, output=-0.846707166504
			11'd1283: out = 32'b10000000000000000110110010100101; // input=-1.013671875, output=-0.848779057547
			11'd1284: out = 32'b10000000000000000110110011101000; // input=-1.017578125, output=-0.850837997266
			11'd1285: out = 32'b10000000000000000110110100101011; // input=-1.021484375, output=-0.852883954244
			11'd1286: out = 32'b10000000000000000110110101101110; // input=-1.025390625, output=-0.854916897262
			11'd1287: out = 32'b10000000000000000110110110110000; // input=-1.029296875, output=-0.8569367953
			11'd1288: out = 32'b10000000000000000110110111110010; // input=-1.033203125, output=-0.858943617537
			11'd1289: out = 32'b10000000000000000110111000110011; // input=-1.037109375, output=-0.860937333352
			11'd1290: out = 32'b10000000000000000110111001110100; // input=-1.041015625, output=-0.862917912321
			11'd1291: out = 32'b10000000000000000110111010110101; // input=-1.044921875, output=-0.864885324225
			11'd1292: out = 32'b10000000000000000110111011110101; // input=-1.048828125, output=-0.866839539044
			11'd1293: out = 32'b10000000000000000110111100110100; // input=-1.052734375, output=-0.868780526957
			11'd1294: out = 32'b10000000000000000110111101110011; // input=-1.056640625, output=-0.870708258348
			11'd1295: out = 32'b10000000000000000110111110110010; // input=-1.060546875, output=-0.872622703803
			11'd1296: out = 32'b10000000000000000110111111110000; // input=-1.064453125, output=-0.874523834109
			11'd1297: out = 32'b10000000000000000111000000101110; // input=-1.068359375, output=-0.876411620257
			11'd1298: out = 32'b10000000000000000111000001101100; // input=-1.072265625, output=-0.878286033441
			11'd1299: out = 32'b10000000000000000111000010101001; // input=-1.076171875, output=-0.880147045062
			11'd1300: out = 32'b10000000000000000111000011100101; // input=-1.080078125, output=-0.881994626722
			11'd1301: out = 32'b10000000000000000111000100100001; // input=-1.083984375, output=-0.883828750229
			11'd1302: out = 32'b10000000000000000111000101011101; // input=-1.087890625, output=-0.885649387596
			11'd1303: out = 32'b10000000000000000111000110011000; // input=-1.091796875, output=-0.887456511044
			11'd1304: out = 32'b10000000000000000111000111010011; // input=-1.095703125, output=-0.889250092997
			11'd1305: out = 32'b10000000000000000111001000001101; // input=-1.099609375, output=-0.891030106087
			11'd1306: out = 32'b10000000000000000111001001000111; // input=-1.103515625, output=-0.892796523155
			11'd1307: out = 32'b10000000000000000111001010000001; // input=-1.107421875, output=-0.894549317246
			11'd1308: out = 32'b10000000000000000111001010111010; // input=-1.111328125, output=-0.896288461615
			11'd1309: out = 32'b10000000000000000111001011110010; // input=-1.115234375, output=-0.898013929725
			11'd1310: out = 32'b10000000000000000111001100101010; // input=-1.119140625, output=-0.899725695247
			11'd1311: out = 32'b10000000000000000111001101100010; // input=-1.123046875, output=-0.901423732062
			11'd1312: out = 32'b10000000000000000111001110011001; // input=-1.126953125, output=-0.90310801426
			11'd1313: out = 32'b10000000000000000111001111010000; // input=-1.130859375, output=-0.90477851614
			11'd1314: out = 32'b10000000000000000111010000000110; // input=-1.134765625, output=-0.906435212214
			11'd1315: out = 32'b10000000000000000111010000111100; // input=-1.138671875, output=-0.908078077202
			11'd1316: out = 32'b10000000000000000111010001110001; // input=-1.142578125, output=-0.909707086035
			11'd1317: out = 32'b10000000000000000111010010100110; // input=-1.146484375, output=-0.911322213858
			11'd1318: out = 32'b10000000000000000111010011011011; // input=-1.150390625, output=-0.912923436025
			11'd1319: out = 32'b10000000000000000111010100001111; // input=-1.154296875, output=-0.914510728103
			11'd1320: out = 32'b10000000000000000111010101000010; // input=-1.158203125, output=-0.916084065873
			11'd1321: out = 32'b10000000000000000111010101110101; // input=-1.162109375, output=-0.917643425327
			11'd1322: out = 32'b10000000000000000111010110101000; // input=-1.166015625, output=-0.919188782671
			11'd1323: out = 32'b10000000000000000111010111011010; // input=-1.169921875, output=-0.920720114326
			11'd1324: out = 32'b10000000000000000111011000001100; // input=-1.173828125, output=-0.922237396924
			11'd1325: out = 32'b10000000000000000111011000111101; // input=-1.177734375, output=-0.923740607315
			11'd1326: out = 32'b10000000000000000111011001101110; // input=-1.181640625, output=-0.92522972256
			11'd1327: out = 32'b10000000000000000111011010011110; // input=-1.185546875, output=-0.926704719938
			11'd1328: out = 32'b10000000000000000111011011001110; // input=-1.189453125, output=-0.928165576942
			11'd1329: out = 32'b10000000000000000111011011111110; // input=-1.193359375, output=-0.929612271281
			11'd1330: out = 32'b10000000000000000111011100101100; // input=-1.197265625, output=-0.931044780881
			11'd1331: out = 32'b10000000000000000111011101011011; // input=-1.201171875, output=-0.932463083883
			11'd1332: out = 32'b10000000000000000111011110001001; // input=-1.205078125, output=-0.933867158646
			11'd1333: out = 32'b10000000000000000111011110110111; // input=-1.208984375, output=-0.935256983744
			11'd1334: out = 32'b10000000000000000111011111100100; // input=-1.212890625, output=-0.936632537972
			11'd1335: out = 32'b10000000000000000111100000010000; // input=-1.216796875, output=-0.93799380034
			11'd1336: out = 32'b10000000000000000111100000111100; // input=-1.220703125, output=-0.939340750076
			11'd1337: out = 32'b10000000000000000111100001101000; // input=-1.224609375, output=-0.940673366629
			11'd1338: out = 32'b10000000000000000111100010010011; // input=-1.228515625, output=-0.941991629663
			11'd1339: out = 32'b10000000000000000111100010111110; // input=-1.232421875, output=-0.943295519063
			11'd1340: out = 32'b10000000000000000111100011101000; // input=-1.236328125, output=-0.944585014935
			11'd1341: out = 32'b10000000000000000111100100010010; // input=-1.240234375, output=-0.945860097601
			11'd1342: out = 32'b10000000000000000111100100111011; // input=-1.244140625, output=-0.947120747606
			11'd1343: out = 32'b10000000000000000111100101100100; // input=-1.248046875, output=-0.948366945714
			11'd1344: out = 32'b10000000000000000111100110001100; // input=-1.251953125, output=-0.949598672909
			11'd1345: out = 32'b10000000000000000111100110110100; // input=-1.255859375, output=-0.950815910397
			11'd1346: out = 32'b10000000000000000111100111011100; // input=-1.259765625, output=-0.952018639603
			11'd1347: out = 32'b10000000000000000111101000000011; // input=-1.263671875, output=-0.953206842177
			11'd1348: out = 32'b10000000000000000111101000101001; // input=-1.267578125, output=-0.954380499987
			11'd1349: out = 32'b10000000000000000111101001001111; // input=-1.271484375, output=-0.955539595124
			11'd1350: out = 32'b10000000000000000111101001110101; // input=-1.275390625, output=-0.956684109903
			11'd1351: out = 32'b10000000000000000111101010011010; // input=-1.279296875, output=-0.95781402686
			11'd1352: out = 32'b10000000000000000111101010111110; // input=-1.283203125, output=-0.958929328753
			11'd1353: out = 32'b10000000000000000111101011100010; // input=-1.287109375, output=-0.960029998564
			11'd1354: out = 32'b10000000000000000111101100000110; // input=-1.291015625, output=-0.961116019499
			11'd1355: out = 32'b10000000000000000111101100101001; // input=-1.294921875, output=-0.962187374985
			11'd1356: out = 32'b10000000000000000111101101001100; // input=-1.298828125, output=-0.963244048676
			11'd1357: out = 32'b10000000000000000111101101101110; // input=-1.302734375, output=-0.964286024448
			11'd1358: out = 32'b10000000000000000111101110001111; // input=-1.306640625, output=-0.965313286402
			11'd1359: out = 32'b10000000000000000111101110110001; // input=-1.310546875, output=-0.966325818863
			11'd1360: out = 32'b10000000000000000111101111010001; // input=-1.314453125, output=-0.96732360638
			11'd1361: out = 32'b10000000000000000111101111110001; // input=-1.318359375, output=-0.96830663373
			11'd1362: out = 32'b10000000000000000111110000010001; // input=-1.322265625, output=-0.969274885911
			11'd1363: out = 32'b10000000000000000111110000110000; // input=-1.326171875, output=-0.970228348151
			11'd1364: out = 32'b10000000000000000111110001001111; // input=-1.330078125, output=-0.971167005899
			11'd1365: out = 32'b10000000000000000111110001101101; // input=-1.333984375, output=-0.972090844834
			11'd1366: out = 32'b10000000000000000111110010001011; // input=-1.337890625, output=-0.972999850858
			11'd1367: out = 32'b10000000000000000111110010101001; // input=-1.341796875, output=-0.973894010102
			11'd1368: out = 32'b10000000000000000111110011000101; // input=-1.345703125, output=-0.974773308922
			11'd1369: out = 32'b10000000000000000111110011100010; // input=-1.349609375, output=-0.9756377339
			11'd1370: out = 32'b10000000000000000111110011111110; // input=-1.353515625, output=-0.976487271847
			11'd1371: out = 32'b10000000000000000111110100011001; // input=-1.357421875, output=-0.977321909799
			11'd1372: out = 32'b10000000000000000111110100110100; // input=-1.361328125, output=-0.978141635021
			11'd1373: out = 32'b10000000000000000111110101001110; // input=-1.365234375, output=-0.978946435006
			11'd1374: out = 32'b10000000000000000111110101101000; // input=-1.369140625, output=-0.979736297472
			11'd1375: out = 32'b10000000000000000111110110000001; // input=-1.373046875, output=-0.980511210368
			11'd1376: out = 32'b10000000000000000111110110011010; // input=-1.376953125, output=-0.981271161869
			11'd1377: out = 32'b10000000000000000111110110110011; // input=-1.380859375, output=-0.98201614038
			11'd1378: out = 32'b10000000000000000111110111001011; // input=-1.384765625, output=-0.982746134532
			11'd1379: out = 32'b10000000000000000111110111100010; // input=-1.388671875, output=-0.983461133188
			11'd1380: out = 32'b10000000000000000111110111111001; // input=-1.392578125, output=-0.984161125436
			11'd1381: out = 32'b10000000000000000111111000001111; // input=-1.396484375, output=-0.984846100597
			11'd1382: out = 32'b10000000000000000111111000100101; // input=-1.400390625, output=-0.985516048218
			11'd1383: out = 32'b10000000000000000111111000111011; // input=-1.404296875, output=-0.986170958077
			11'd1384: out = 32'b10000000000000000111111001010000; // input=-1.408203125, output=-0.98681082018
			11'd1385: out = 32'b10000000000000000111111001100100; // input=-1.412109375, output=-0.987435624764
			11'd1386: out = 32'b10000000000000000111111001111000; // input=-1.416015625, output=-0.988045362295
			11'd1387: out = 32'b10000000000000000111111010001100; // input=-1.419921875, output=-0.98864002347
			11'd1388: out = 32'b10000000000000000111111010011111; // input=-1.423828125, output=-0.989219599214
			11'd1389: out = 32'b10000000000000000111111010110001; // input=-1.427734375, output=-0.989784080684
			11'd1390: out = 32'b10000000000000000111111011000011; // input=-1.431640625, output=-0.990333459267
			11'd1391: out = 32'b10000000000000000111111011010101; // input=-1.435546875, output=-0.99086772658
			11'd1392: out = 32'b10000000000000000111111011100110; // input=-1.439453125, output=-0.991386874471
			11'd1393: out = 32'b10000000000000000111111011110110; // input=-1.443359375, output=-0.991890895017
			11'd1394: out = 32'b10000000000000000111111100000110; // input=-1.447265625, output=-0.992379780529
			11'd1395: out = 32'b10000000000000000111111100010110; // input=-1.451171875, output=-0.992853523546
			11'd1396: out = 32'b10000000000000000111111100100101; // input=-1.455078125, output=-0.99331211684
			11'd1397: out = 32'b10000000000000000111111100110011; // input=-1.458984375, output=-0.993755553414
			11'd1398: out = 32'b10000000000000000111111101000001; // input=-1.462890625, output=-0.9941838265
			11'd1399: out = 32'b10000000000000000111111101001111; // input=-1.466796875, output=-0.994596929564
			11'd1400: out = 32'b10000000000000000111111101011100; // input=-1.470703125, output=-0.994994856303
			11'd1401: out = 32'b10000000000000000111111101101001; // input=-1.474609375, output=-0.995377600644
			11'd1402: out = 32'b10000000000000000111111101110101; // input=-1.478515625, output=-0.995745156748
			11'd1403: out = 32'b10000000000000000111111110000000; // input=-1.482421875, output=-0.996097519006
			11'd1404: out = 32'b10000000000000000111111110001011; // input=-1.486328125, output=-0.996434682041
			11'd1405: out = 32'b10000000000000000111111110010110; // input=-1.490234375, output=-0.996756640709
			11'd1406: out = 32'b10000000000000000111111110100000; // input=-1.494140625, output=-0.997063390097
			11'd1407: out = 32'b10000000000000000111111110101001; // input=-1.498046875, output=-0.997354925525
			11'd1408: out = 32'b10000000000000000111111110110010; // input=-1.501953125, output=-0.997631242543
			11'd1409: out = 32'b10000000000000000111111110111011; // input=-1.505859375, output=-0.997892336936
			11'd1410: out = 32'b10000000000000000111111111000011; // input=-1.509765625, output=-0.99813820472
			11'd1411: out = 32'b10000000000000000111111111001011; // input=-1.513671875, output=-0.998368842143
			11'd1412: out = 32'b10000000000000000111111111010010; // input=-1.517578125, output=-0.998584245685
			11'd1413: out = 32'b10000000000000000111111111011000; // input=-1.521484375, output=-0.998784412061
			11'd1414: out = 32'b10000000000000000111111111011110; // input=-1.525390625, output=-0.998969338215
			11'd1415: out = 32'b10000000000000000111111111100100; // input=-1.529296875, output=-0.999139021326
			11'd1416: out = 32'b10000000000000000111111111101001; // input=-1.533203125, output=-0.999293458805
			11'd1417: out = 32'b10000000000000000111111111101101; // input=-1.537109375, output=-0.999432648295
			11'd1418: out = 32'b10000000000000000111111111110001; // input=-1.541015625, output=-0.999556587673
			11'd1419: out = 32'b10000000000000000111111111110101; // input=-1.544921875, output=-0.999665275047
			11'd1420: out = 32'b10000000000000000111111111111000; // input=-1.548828125, output=-0.999758708759
			11'd1421: out = 32'b10000000000000000111111111111011; // input=-1.552734375, output=-0.999836887383
			11'd1422: out = 32'b10000000000000000111111111111101; // input=-1.556640625, output=-0.999899809726
			11'd1423: out = 32'b10000000000000000111111111111110; // input=-1.560546875, output=-0.999947474829
			11'd1424: out = 32'b10000000000000000111111111111111; // input=-1.564453125, output=-0.999979881963
			11'd1425: out = 32'b10000000000000000111111111111111; // input=-1.568359375, output=-0.999997030634
			11'd1426: out = 32'b10000000000000000111111111111111; // input=-1.572265625, output=-0.999998920582
			11'd1427: out = 32'b10000000000000000111111111111111; // input=-1.576171875, output=-0.999985551776
			11'd1428: out = 32'b10000000000000000111111111111111; // input=-1.580078125, output=-0.99995692442
			11'd1429: out = 32'b10000000000000000111111111111101; // input=-1.583984375, output=-0.999913038953
			11'd1430: out = 32'b10000000000000000111111111111011; // input=-1.587890625, output=-0.999853896042
			11'd1431: out = 32'b10000000000000000111111111111001; // input=-1.591796875, output=-0.999779496592
			11'd1432: out = 32'b10000000000000000111111111110110; // input=-1.595703125, output=-0.999689841736
			11'd1433: out = 32'b10000000000000000111111111110010; // input=-1.599609375, output=-0.999584932843
			11'd1434: out = 32'b10000000000000000111111111101110; // input=-1.603515625, output=-0.999464771514
			11'd1435: out = 32'b10000000000000000111111111101010; // input=-1.607421875, output=-0.999329359583
			11'd1436: out = 32'b10000000000000000111111111100101; // input=-1.611328125, output=-0.999178699114
			11'd1437: out = 32'b10000000000000000111111111100000; // input=-1.615234375, output=-0.999012792408
			11'd1438: out = 32'b10000000000000000111111111011010; // input=-1.619140625, output=-0.998831641997
			11'd1439: out = 32'b10000000000000000111111111010011; // input=-1.623046875, output=-0.998635250643
			11'd1440: out = 32'b10000000000000000111111111001100; // input=-1.626953125, output=-0.998423621343
			11'd1441: out = 32'b10000000000000000111111111000101; // input=-1.630859375, output=-0.998196757328
			11'd1442: out = 32'b10000000000000000111111110111101; // input=-1.634765625, output=-0.997954662059
			11'd1443: out = 32'b10000000000000000111111110110101; // input=-1.638671875, output=-0.997697339229
			11'd1444: out = 32'b10000000000000000111111110101100; // input=-1.642578125, output=-0.997424792765
			11'd1445: out = 32'b10000000000000000111111110100010; // input=-1.646484375, output=-0.997137026826
			11'd1446: out = 32'b10000000000000000111111110011000; // input=-1.650390625, output=-0.996834045803
			11'd1447: out = 32'b10000000000000000111111110001110; // input=-1.654296875, output=-0.996515854318
			11'd1448: out = 32'b10000000000000000111111110000011; // input=-1.658203125, output=-0.996182457228
			11'd1449: out = 32'b10000000000000000111111101110111; // input=-1.662109375, output=-0.995833859619
			11'd1450: out = 32'b10000000000000000111111101101100; // input=-1.666015625, output=-0.995470066811
			11'd1451: out = 32'b10000000000000000111111101011111; // input=-1.669921875, output=-0.995091084354
			11'd1452: out = 32'b10000000000000000111111101010010; // input=-1.673828125, output=-0.994696918032
			11'd1453: out = 32'b10000000000000000111111101000101; // input=-1.677734375, output=-0.994287573858
			11'd1454: out = 32'b10000000000000000111111100110111; // input=-1.681640625, output=-0.99386305808
			11'd1455: out = 32'b10000000000000000111111100101000; // input=-1.685546875, output=-0.993423377174
			11'd1456: out = 32'b10000000000000000111111100011010; // input=-1.689453125, output=-0.992968537849
			11'd1457: out = 32'b10000000000000000111111100001010; // input=-1.693359375, output=-0.992498547046
			11'd1458: out = 32'b10000000000000000111111011111010; // input=-1.697265625, output=-0.992013411937
			11'd1459: out = 32'b10000000000000000111111011101010; // input=-1.701171875, output=-0.991513139923
			11'd1460: out = 32'b10000000000000000111111011011001; // input=-1.705078125, output=-0.990997738639
			11'd1461: out = 32'b10000000000000000111111011001000; // input=-1.708984375, output=-0.990467215948
			11'd1462: out = 32'b10000000000000000111111010110110; // input=-1.712890625, output=-0.989921579947
			11'd1463: out = 32'b10000000000000000111111010100011; // input=-1.716796875, output=-0.98936083896
			11'd1464: out = 32'b10000000000000000111111010010001; // input=-1.720703125, output=-0.988785001544
			11'd1465: out = 32'b10000000000000000111111001111101; // input=-1.724609375, output=-0.988194076485
			11'd1466: out = 32'b10000000000000000111111001101001; // input=-1.728515625, output=-0.9875880728
			11'd1467: out = 32'b10000000000000000111111001010101; // input=-1.732421875, output=-0.986966999737
			11'd1468: out = 32'b10000000000000000111111001000000; // input=-1.736328125, output=-0.986330866772
			11'd1469: out = 32'b10000000000000000111111000101011; // input=-1.740234375, output=-0.98567968361
			11'd1470: out = 32'b10000000000000000111111000010101; // input=-1.744140625, output=-0.98501346019
			11'd1471: out = 32'b10000000000000000111110111111111; // input=-1.748046875, output=-0.984332206676
			11'd1472: out = 32'b10000000000000000111110111101000; // input=-1.751953125, output=-0.983635933464
			11'd1473: out = 32'b10000000000000000111110111010000; // input=-1.755859375, output=-0.982924651178
			11'd1474: out = 32'b10000000000000000111110110111001; // input=-1.759765625, output=-0.982198370671
			11'd1475: out = 32'b10000000000000000111110110100000; // input=-1.763671875, output=-0.981457103025
			11'd1476: out = 32'b10000000000000000111110110001000; // input=-1.767578125, output=-0.980700859551
			11'd1477: out = 32'b10000000000000000111110101101110; // input=-1.771484375, output=-0.979929651789
			11'd1478: out = 32'b10000000000000000111110101010101; // input=-1.775390625, output=-0.979143491506
			11'd1479: out = 32'b10000000000000000111110100111010; // input=-1.779296875, output=-0.978342390698
			11'd1480: out = 32'b10000000000000000111110100100000; // input=-1.783203125, output=-0.977526361588
			11'd1481: out = 32'b10000000000000000111110100000100; // input=-1.787109375, output=-0.976695416629
			11'd1482: out = 32'b10000000000000000111110011101001; // input=-1.791015625, output=-0.9758495685
			11'd1483: out = 32'b10000000000000000111110011001100; // input=-1.794921875, output=-0.974988830107
			11'd1484: out = 32'b10000000000000000111110010110000; // input=-1.798828125, output=-0.974113214584
			11'd1485: out = 32'b10000000000000000111110010010011; // input=-1.802734375, output=-0.973222735292
			11'd1486: out = 32'b10000000000000000111110001110101; // input=-1.806640625, output=-0.972317405818
			11'd1487: out = 32'b10000000000000000111110001010111; // input=-1.810546875, output=-0.971397239977
			11'd1488: out = 32'b10000000000000000111110000111000; // input=-1.814453125, output=-0.970462251809
			11'd1489: out = 32'b10000000000000000111110000011001; // input=-1.818359375, output=-0.969512455581
			11'd1490: out = 32'b10000000000000000111101111111001; // input=-1.822265625, output=-0.968547865786
			11'd1491: out = 32'b10000000000000000111101111011001; // input=-1.826171875, output=-0.967568497142
			11'd1492: out = 32'b10000000000000000111101110111001; // input=-1.830078125, output=-0.966574364594
			11'd1493: out = 32'b10000000000000000111101110011000; // input=-1.833984375, output=-0.96556548331
			11'd1494: out = 32'b10000000000000000111101101110110; // input=-1.837890625, output=-0.964541868684
			11'd1495: out = 32'b10000000000000000111101101010100; // input=-1.841796875, output=-0.963503536336
			11'd1496: out = 32'b10000000000000000111101100110010; // input=-1.845703125, output=-0.96245050211
			11'd1497: out = 32'b10000000000000000111101100001111; // input=-1.849609375, output=-0.961382782073
			11'd1498: out = 32'b10000000000000000111101011101011; // input=-1.853515625, output=-0.960300392518
			11'd1499: out = 32'b10000000000000000111101011000111; // input=-1.857421875, output=-0.95920334996
			11'd1500: out = 32'b10000000000000000111101010100011; // input=-1.861328125, output=-0.95809167114
			11'd1501: out = 32'b10000000000000000111101001111110; // input=-1.865234375, output=-0.956965373019
			11'd1502: out = 32'b10000000000000000111101001011000; // input=-1.869140625, output=-0.955824472784
			11'd1503: out = 32'b10000000000000000111101000110011; // input=-1.873046875, output=-0.954668987843
			11'd1504: out = 32'b10000000000000000111101000001100; // input=-1.876953125, output=-0.953498935829
			11'd1505: out = 32'b10000000000000000111100111100101; // input=-1.880859375, output=-0.952314334593
			11'd1506: out = 32'b10000000000000000111100110111110; // input=-1.884765625, output=-0.951115202213
			11'd1507: out = 32'b10000000000000000111100110010110; // input=-1.888671875, output=-0.949901556985
			11'd1508: out = 32'b10000000000000000111100101101110; // input=-1.892578125, output=-0.948673417428
			11'd1509: out = 32'b10000000000000000111100101000101; // input=-1.896484375, output=-0.947430802281
			11'd1510: out = 32'b10000000000000000111100100011100; // input=-1.900390625, output=-0.946173730507
			11'd1511: out = 32'b10000000000000000111100011110011; // input=-1.904296875, output=-0.944902221285
			11'd1512: out = 32'b10000000000000000111100011001000; // input=-1.908203125, output=-0.943616294018
			11'd1513: out = 32'b10000000000000000111100010011110; // input=-1.912109375, output=-0.942315968327
			11'd1514: out = 32'b10000000000000000111100001110011; // input=-1.916015625, output=-0.941001264054
			11'd1515: out = 32'b10000000000000000111100001000111; // input=-1.919921875, output=-0.939672201259
			11'd1516: out = 32'b10000000000000000111100000011011; // input=-1.923828125, output=-0.938328800223
			11'd1517: out = 32'b10000000000000000111011111101111; // input=-1.927734375, output=-0.936971081444
			11'd1518: out = 32'b10000000000000000111011111000010; // input=-1.931640625, output=-0.935599065638
			11'd1519: out = 32'b10000000000000000111011110010100; // input=-1.935546875, output=-0.934212773742
			11'd1520: out = 32'b10000000000000000111011101100110; // input=-1.939453125, output=-0.932812226909
			11'd1521: out = 32'b10000000000000000111011100111000; // input=-1.943359375, output=-0.931397446509
			11'd1522: out = 32'b10000000000000000111011100001001; // input=-1.947265625, output=-0.929968454129
			11'd1523: out = 32'b10000000000000000111011011011010; // input=-1.951171875, output=-0.928525271575
			11'd1524: out = 32'b10000000000000000111011010101010; // input=-1.955078125, output=-0.927067920868
			11'd1525: out = 32'b10000000000000000111011001111010; // input=-1.958984375, output=-0.925596424245
			11'd1526: out = 32'b10000000000000000111011001001001; // input=-1.962890625, output=-0.92411080416
			11'd1527: out = 32'b10000000000000000111011000011000; // input=-1.966796875, output=-0.92261108328
			11'd1528: out = 32'b10000000000000000111010111100111; // input=-1.970703125, output=-0.921097284491
			11'd1529: out = 32'b10000000000000000111010110110100; // input=-1.974609375, output=-0.91956943089
			11'd1530: out = 32'b10000000000000000111010110000010; // input=-1.978515625, output=-0.918027545791
			11'd1531: out = 32'b10000000000000000111010101001111; // input=-1.982421875, output=-0.916471652721
			11'd1532: out = 32'b10000000000000000111010100011100; // input=-1.986328125, output=-0.914901775422
			11'd1533: out = 32'b10000000000000000111010011101000; // input=-1.990234375, output=-0.913317937847
			11'd1534: out = 32'b10000000000000000111010010110011; // input=-1.994140625, output=-0.911720164164
			11'd1535: out = 32'b10000000000000000111010001111110; // input=-1.998046875, output=-0.910108478752
			11'd1536: out = 32'b10000000000000000111010001001001; // input=-2.001953125, output=-0.908482906206
			11'd1537: out = 32'b10000000000000000111010000010011; // input=-2.005859375, output=-0.906843471327
			11'd1538: out = 32'b10000000000000000111001111011101; // input=-2.009765625, output=-0.905190199134
			11'd1539: out = 32'b10000000000000000111001110100111; // input=-2.013671875, output=-0.903523114851
			11'd1540: out = 32'b10000000000000000111001101110000; // input=-2.017578125, output=-0.901842243918
			11'd1541: out = 32'b10000000000000000111001100111000; // input=-2.021484375, output=-0.900147611981
			11'd1542: out = 32'b10000000000000000111001100000000; // input=-2.025390625, output=-0.898439244899
			11'd1543: out = 32'b10000000000000000111001011001000; // input=-2.029296875, output=-0.89671716874
			11'd1544: out = 32'b10000000000000000111001010001111; // input=-2.033203125, output=-0.89498140978
			11'd1545: out = 32'b10000000000000000111001001010101; // input=-2.037109375, output=-0.893231994505
			11'd1546: out = 32'b10000000000000000111001000011100; // input=-2.041015625, output=-0.891468949608
			11'd1547: out = 32'b10000000000000000111000111100001; // input=-2.044921875, output=-0.889692301992
			11'd1548: out = 32'b10000000000000000111000110100111; // input=-2.048828125, output=-0.887902078767
			11'd1549: out = 32'b10000000000000000111000101101100; // input=-2.052734375, output=-0.886098307248
			11'd1550: out = 32'b10000000000000000111000100110000; // input=-2.056640625, output=-0.884281014959
			11'd1551: out = 32'b10000000000000000111000011110100; // input=-2.060546875, output=-0.882450229629
			11'd1552: out = 32'b10000000000000000111000010111000; // input=-2.064453125, output=-0.880605979195
			11'd1553: out = 32'b10000000000000000111000001111011; // input=-2.068359375, output=-0.878748291797
			11'd1554: out = 32'b10000000000000000111000000111110; // input=-2.072265625, output=-0.876877195782
			11'd1555: out = 32'b10000000000000000111000000000000; // input=-2.076171875, output=-0.874992719699
			11'd1556: out = 32'b10000000000000000110111111000010; // input=-2.080078125, output=-0.873094892304
			11'd1557: out = 32'b10000000000000000110111110000011; // input=-2.083984375, output=-0.871183742555
			11'd1558: out = 32'b10000000000000000110111101000100; // input=-2.087890625, output=-0.869259299614
			11'd1559: out = 32'b10000000000000000110111100000100; // input=-2.091796875, output=-0.867321592845
			11'd1560: out = 32'b10000000000000000110111011000100; // input=-2.095703125, output=-0.865370651816
			11'd1561: out = 32'b10000000000000000110111010000100; // input=-2.099609375, output=-0.863406506296
			11'd1562: out = 32'b10000000000000000110111001000011; // input=-2.103515625, output=-0.861429186254
			11'd1563: out = 32'b10000000000000000110111000000010; // input=-2.107421875, output=-0.859438721864
			11'd1564: out = 32'b10000000000000000110110111000000; // input=-2.111328125, output=-0.857435143495
			11'd1565: out = 32'b10000000000000000110110101111110; // input=-2.115234375, output=-0.855418481721
			11'd1566: out = 32'b10000000000000000110110100111100; // input=-2.119140625, output=-0.853388767314
			11'd1567: out = 32'b10000000000000000110110011111001; // input=-2.123046875, output=-0.851346031244
			11'd1568: out = 32'b10000000000000000110110010110110; // input=-2.126953125, output=-0.849290304681
			11'd1569: out = 32'b10000000000000000110110001110010; // input=-2.130859375, output=-0.847221618993
			11'd1570: out = 32'b10000000000000000110110000101110; // input=-2.134765625, output=-0.845140005746
			11'd1571: out = 32'b10000000000000000110101111101001; // input=-2.138671875, output=-0.843045496701
			11'd1572: out = 32'b10000000000000000110101110100100; // input=-2.142578125, output=-0.84093812382
			11'd1573: out = 32'b10000000000000000110101101011110; // input=-2.146484375, output=-0.838817919257
			11'd1574: out = 32'b10000000000000000110101100011000; // input=-2.150390625, output=-0.836684915366
			11'd1575: out = 32'b10000000000000000110101011010010; // input=-2.154296875, output=-0.834539144691
			11'd1576: out = 32'b10000000000000000110101010001011; // input=-2.158203125, output=-0.832380639976
			11'd1577: out = 32'b10000000000000000110101001000100; // input=-2.162109375, output=-0.830209434157
			11'd1578: out = 32'b10000000000000000110100111111101; // input=-2.166015625, output=-0.828025560363
			11'd1579: out = 32'b10000000000000000110100110110101; // input=-2.169921875, output=-0.825829051918
			11'd1580: out = 32'b10000000000000000110100101101100; // input=-2.173828125, output=-0.823619942338
			11'd1581: out = 32'b10000000000000000110100100100100; // input=-2.177734375, output=-0.82139826533
			11'd1582: out = 32'b10000000000000000110100011011010; // input=-2.181640625, output=-0.819164054796
			11'd1583: out = 32'b10000000000000000110100010010001; // input=-2.185546875, output=-0.816917344826
			11'd1584: out = 32'b10000000000000000110100001000111; // input=-2.189453125, output=-0.814658169702
			11'd1585: out = 32'b10000000000000000110011111111100; // input=-2.193359375, output=-0.812386563897
			11'd1586: out = 32'b10000000000000000110011110110001; // input=-2.197265625, output=-0.810102562073
			11'd1587: out = 32'b10000000000000000110011101100110; // input=-2.201171875, output=-0.80780619908
			11'd1588: out = 32'b10000000000000000110011100011011; // input=-2.205078125, output=-0.805497509959
			11'd1589: out = 32'b10000000000000000110011011001110; // input=-2.208984375, output=-0.803176529936
			11'd1590: out = 32'b10000000000000000110011010000010; // input=-2.212890625, output=-0.800843294428
			11'd1591: out = 32'b10000000000000000110011000110101; // input=-2.216796875, output=-0.798497839037
			11'd1592: out = 32'b10000000000000000110010111101000; // input=-2.220703125, output=-0.796140199551
			11'd1593: out = 32'b10000000000000000110010110011010; // input=-2.224609375, output=-0.793770411945
			11'd1594: out = 32'b10000000000000000110010101001100; // input=-2.228515625, output=-0.791388512379
			11'd1595: out = 32'b10000000000000000110010011111110; // input=-2.232421875, output=-0.788994537198
			11'd1596: out = 32'b10000000000000000110010010101111; // input=-2.236328125, output=-0.786588522931
			11'd1597: out = 32'b10000000000000000110010001100000; // input=-2.240234375, output=-0.784170506291
			11'd1598: out = 32'b10000000000000000110010000010000; // input=-2.244140625, output=-0.781740524174
			11'd1599: out = 32'b10000000000000000110001111000000; // input=-2.248046875, output=-0.779298613658
			11'd1600: out = 32'b10000000000000000110001101110000; // input=-2.251953125, output=-0.776844812005
			11'd1601: out = 32'b10000000000000000110001100011111; // input=-2.255859375, output=-0.774379156655
			11'd1602: out = 32'b10000000000000000110001011001110; // input=-2.259765625, output=-0.771901685232
			11'd1603: out = 32'b10000000000000000110001001111100; // input=-2.263671875, output=-0.769412435539
			11'd1604: out = 32'b10000000000000000110001000101010; // input=-2.267578125, output=-0.766911445559
			11'd1605: out = 32'b10000000000000000110000111011000; // input=-2.271484375, output=-0.764398753454
			11'd1606: out = 32'b10000000000000000110000110000101; // input=-2.275390625, output=-0.761874397564
			11'd1607: out = 32'b10000000000000000110000100110010; // input=-2.279296875, output=-0.759338416409
			11'd1608: out = 32'b10000000000000000110000011011111; // input=-2.283203125, output=-0.756790848683
			11'd1609: out = 32'b10000000000000000110000010001011; // input=-2.287109375, output=-0.75423173326
			11'd1610: out = 32'b10000000000000000110000000110110; // input=-2.291015625, output=-0.751661109189
			11'd1611: out = 32'b10000000000000000101111111100010; // input=-2.294921875, output=-0.749079015694
			11'd1612: out = 32'b10000000000000000101111110001101; // input=-2.298828125, output=-0.746485492175
			11'd1613: out = 32'b10000000000000000101111100110111; // input=-2.302734375, output=-0.743880578206
			11'd1614: out = 32'b10000000000000000101111011100010; // input=-2.306640625, output=-0.741264313535
			11'd1615: out = 32'b10000000000000000101111010001100; // input=-2.310546875, output=-0.738636738082
			11'd1616: out = 32'b10000000000000000101111000110101; // input=-2.314453125, output=-0.735997891941
			11'd1617: out = 32'b10000000000000000101110111011110; // input=-2.318359375, output=-0.733347815378
			11'd1618: out = 32'b10000000000000000101110110000111; // input=-2.322265625, output=-0.730686548829
			11'd1619: out = 32'b10000000000000000101110100110000; // input=-2.326171875, output=-0.728014132903
			11'd1620: out = 32'b10000000000000000101110011011000; // input=-2.330078125, output=-0.725330608377
			11'd1621: out = 32'b10000000000000000101110001111111; // input=-2.333984375, output=-0.722636016198
			11'd1622: out = 32'b10000000000000000101110000100111; // input=-2.337890625, output=-0.719930397482
			11'd1623: out = 32'b10000000000000000101101111001110; // input=-2.341796875, output=-0.717213793515
			11'd1624: out = 32'b10000000000000000101101101110100; // input=-2.345703125, output=-0.714486245747
			11'd1625: out = 32'b10000000000000000101101100011011; // input=-2.349609375, output=-0.711747795798
			11'd1626: out = 32'b10000000000000000101101011000000; // input=-2.353515625, output=-0.708998485454
			11'd1627: out = 32'b10000000000000000101101001100110; // input=-2.357421875, output=-0.706238356665
			11'd1628: out = 32'b10000000000000000101101000001011; // input=-2.361328125, output=-0.703467451548
			11'd1629: out = 32'b10000000000000000101100110110000; // input=-2.365234375, output=-0.700685812383
			11'd1630: out = 32'b10000000000000000101100101010101; // input=-2.369140625, output=-0.697893481614
			11'd1631: out = 32'b10000000000000000101100011111001; // input=-2.373046875, output=-0.69509050185
			11'd1632: out = 32'b10000000000000000101100010011101; // input=-2.376953125, output=-0.692276915859
			11'd1633: out = 32'b10000000000000000101100001000000; // input=-2.380859375, output=-0.689452766575
			11'd1634: out = 32'b10000000000000000101011111100011; // input=-2.384765625, output=-0.68661809709
			11'd1635: out = 32'b10000000000000000101011110000110; // input=-2.388671875, output=-0.683772950657
			11'd1636: out = 32'b10000000000000000101011100101000; // input=-2.392578125, output=-0.680917370691
			11'd1637: out = 32'b10000000000000000101011011001010; // input=-2.396484375, output=-0.678051400763
			11'd1638: out = 32'b10000000000000000101011001101100; // input=-2.400390625, output=-0.675175084605
			11'd1639: out = 32'b10000000000000000101011000001110; // input=-2.404296875, output=-0.672288466105
			11'd1640: out = 32'b10000000000000000101010110101111; // input=-2.408203125, output=-0.669391589311
			11'd1641: out = 32'b10000000000000000101010101001111; // input=-2.412109375, output=-0.666484498425
			11'd1642: out = 32'b10000000000000000101010011110000; // input=-2.416015625, output=-0.663567237806
			11'd1643: out = 32'b10000000000000000101010010010000; // input=-2.419921875, output=-0.660639851967
			11'd1644: out = 32'b10000000000000000101010000110000; // input=-2.423828125, output=-0.657702385576
			11'd1645: out = 32'b10000000000000000101001111001111; // input=-2.427734375, output=-0.654754883457
			11'd1646: out = 32'b10000000000000000101001101101110; // input=-2.431640625, output=-0.651797390583
			11'd1647: out = 32'b10000000000000000101001100001101; // input=-2.435546875, output=-0.648829952083
			11'd1648: out = 32'b10000000000000000101001010101011; // input=-2.439453125, output=-0.645852613236
			11'd1649: out = 32'b10000000000000000101001001001001; // input=-2.443359375, output=-0.642865419473
			11'd1650: out = 32'b10000000000000000101000111100111; // input=-2.447265625, output=-0.639868416375
			11'd1651: out = 32'b10000000000000000101000110000101; // input=-2.451171875, output=-0.636861649672
			11'd1652: out = 32'b10000000000000000101000100100010; // input=-2.455078125, output=-0.633845165244
			11'd1653: out = 32'b10000000000000000101000010111111; // input=-2.458984375, output=-0.630819009118
			11'd1654: out = 32'b10000000000000000101000001011011; // input=-2.462890625, output=-0.62778322747
			11'd1655: out = 32'b10000000000000000100111111110111; // input=-2.466796875, output=-0.624737866623
			11'd1656: out = 32'b10000000000000000100111110010011; // input=-2.470703125, output=-0.621682973045
			11'd1657: out = 32'b10000000000000000100111100101111; // input=-2.474609375, output=-0.618618593349
			11'd1658: out = 32'b10000000000000000100111011001010; // input=-2.478515625, output=-0.615544774295
			11'd1659: out = 32'b10000000000000000100111001100101; // input=-2.482421875, output=-0.612461562784
			11'd1660: out = 32'b10000000000000000100111000000000; // input=-2.486328125, output=-0.609369005864
			11'd1661: out = 32'b10000000000000000100110110011010; // input=-2.490234375, output=-0.606267150722
			11'd1662: out = 32'b10000000000000000100110100110100; // input=-2.494140625, output=-0.60315604469
			11'd1663: out = 32'b10000000000000000100110011001110; // input=-2.498046875, output=-0.600035735239
			11'd1664: out = 32'b10000000000000000100110001100111; // input=-2.501953125, output=-0.59690626998
			11'd1665: out = 32'b10000000000000000100110000000001; // input=-2.505859375, output=-0.593767696666
			11'd1666: out = 32'b10000000000000000100101110011001; // input=-2.509765625, output=-0.590620063188
			11'd1667: out = 32'b10000000000000000100101100110010; // input=-2.513671875, output=-0.587463417574
			11'd1668: out = 32'b10000000000000000100101011001010; // input=-2.517578125, output=-0.584297807991
			11'd1669: out = 32'b10000000000000000100101001100010; // input=-2.521484375, output=-0.581123282743
			11'd1670: out = 32'b10000000000000000100100111111010; // input=-2.525390625, output=-0.577939890268
			11'd1671: out = 32'b10000000000000000100100110010001; // input=-2.529296875, output=-0.574747679141
			11'd1672: out = 32'b10000000000000000100100100101000; // input=-2.533203125, output=-0.571546698072
			11'd1673: out = 32'b10000000000000000100100010111111; // input=-2.537109375, output=-0.568336995904
			11'd1674: out = 32'b10000000000000000100100001010110; // input=-2.541015625, output=-0.565118621612
			11'd1675: out = 32'b10000000000000000100011111101100; // input=-2.544921875, output=-0.561891624306
			11'd1676: out = 32'b10000000000000000100011110000010; // input=-2.548828125, output=-0.558656053224
			11'd1677: out = 32'b10000000000000000100011100011000; // input=-2.552734375, output=-0.555411957739
			11'd1678: out = 32'b10000000000000000100011010101101; // input=-2.556640625, output=-0.55215938735
			11'd1679: out = 32'b10000000000000000100011001000010; // input=-2.560546875, output=-0.548898391689
			11'd1680: out = 32'b10000000000000000100010111010111; // input=-2.564453125, output=-0.545629020513
			11'd1681: out = 32'b10000000000000000100010101101100; // input=-2.568359375, output=-0.54235132371
			11'd1682: out = 32'b10000000000000000100010100000000; // input=-2.572265625, output=-0.539065351293
			11'd1683: out = 32'b10000000000000000100010010010100; // input=-2.576171875, output=-0.535771153402
			11'd1684: out = 32'b10000000000000000100010000101000; // input=-2.580078125, output=-0.532468780302
			11'd1685: out = 32'b10000000000000000100001110111011; // input=-2.583984375, output=-0.529158282384
			11'd1686: out = 32'b10000000000000000100001101001111; // input=-2.587890625, output=-0.525839710162
			11'd1687: out = 32'b10000000000000000100001011100010; // input=-2.591796875, output=-0.522513114272
			11'd1688: out = 32'b10000000000000000100001001110100; // input=-2.595703125, output=-0.519178545475
			11'd1689: out = 32'b10000000000000000100001000000111; // input=-2.599609375, output=-0.515836054653
			11'd1690: out = 32'b10000000000000000100000110011001; // input=-2.603515625, output=-0.512485692806
			11'd1691: out = 32'b10000000000000000100000100101011; // input=-2.607421875, output=-0.509127511059
			11'd1692: out = 32'b10000000000000000100000010111101; // input=-2.611328125, output=-0.505761560652
			11'd1693: out = 32'b10000000000000000100000001001110; // input=-2.615234375, output=-0.502387892946
			11'd1694: out = 32'b10000000000000000011111111011111; // input=-2.619140625, output=-0.499006559419
			11'd1695: out = 32'b10000000000000000011111101110000; // input=-2.623046875, output=-0.495617611666
			11'd1696: out = 32'b10000000000000000011111100000001; // input=-2.626953125, output=-0.492221101398
			11'd1697: out = 32'b10000000000000000011111010010010; // input=-2.630859375, output=-0.488817080442
			11'd1698: out = 32'b10000000000000000011111000100010; // input=-2.634765625, output=-0.485405600738
			11'd1699: out = 32'b10000000000000000011110110110010; // input=-2.638671875, output=-0.481986714342
			11'd1700: out = 32'b10000000000000000011110101000001; // input=-2.642578125, output=-0.478560473421
			11'd1701: out = 32'b10000000000000000011110011010001; // input=-2.646484375, output=-0.475126930257
			11'd1702: out = 32'b10000000000000000011110001100000; // input=-2.650390625, output=-0.47168613724
			11'd1703: out = 32'b10000000000000000011101111101111; // input=-2.654296875, output=-0.468238146873
			11'd1704: out = 32'b10000000000000000011101101111110; // input=-2.658203125, output=-0.464783011769
			11'd1705: out = 32'b10000000000000000011101100001101; // input=-2.662109375, output=-0.461320784647
			11'd1706: out = 32'b10000000000000000011101010011011; // input=-2.666015625, output=-0.457851518337
			11'd1707: out = 32'b10000000000000000011101000101001; // input=-2.669921875, output=-0.454375265777
			11'd1708: out = 32'b10000000000000000011100110110111; // input=-2.673828125, output=-0.450892080009
			11'd1709: out = 32'b10000000000000000011100101000100; // input=-2.677734375, output=-0.447402014183
			11'd1710: out = 32'b10000000000000000011100011010010; // input=-2.681640625, output=-0.443905121553
			11'd1711: out = 32'b10000000000000000011100001011111; // input=-2.685546875, output=-0.440401455476
			11'd1712: out = 32'b10000000000000000011011111101100; // input=-2.689453125, output=-0.436891069416
			11'd1713: out = 32'b10000000000000000011011101111001; // input=-2.693359375, output=-0.433374016935
			11'd1714: out = 32'b10000000000000000011011100000101; // input=-2.697265625, output=-0.429850351699
			11'd1715: out = 32'b10000000000000000011011010010010; // input=-2.701171875, output=-0.426320127476
			11'd1716: out = 32'b10000000000000000011011000011110; // input=-2.705078125, output=-0.422783398133
			11'd1717: out = 32'b10000000000000000011010110101010; // input=-2.708984375, output=-0.419240217635
			11'd1718: out = 32'b10000000000000000011010100110101; // input=-2.712890625, output=-0.415690640047
			11'd1719: out = 32'b10000000000000000011010011000001; // input=-2.716796875, output=-0.412134719532
			11'd1720: out = 32'b10000000000000000011010001001100; // input=-2.720703125, output=-0.408572510347
			11'd1721: out = 32'b10000000000000000011001111010111; // input=-2.724609375, output=-0.405004066849
			11'd1722: out = 32'b10000000000000000011001101100010; // input=-2.728515625, output=-0.401429443487
			11'd1723: out = 32'b10000000000000000011001011101101; // input=-2.732421875, output=-0.397848694806
			11'd1724: out = 32'b10000000000000000011001001110111; // input=-2.736328125, output=-0.394261875443
			11'd1725: out = 32'b10000000000000000011001000000001; // input=-2.740234375, output=-0.390669040129
			11'd1726: out = 32'b10000000000000000011000110001100; // input=-2.744140625, output=-0.387070243686
			11'd1727: out = 32'b10000000000000000011000100010101; // input=-2.748046875, output=-0.383465541027
			11'd1728: out = 32'b10000000000000000011000010011111; // input=-2.751953125, output=-0.379854987156
			11'd1729: out = 32'b10000000000000000011000000101001; // input=-2.755859375, output=-0.376238637166
			11'd1730: out = 32'b10000000000000000010111110110010; // input=-2.759765625, output=-0.372616546236
			11'd1731: out = 32'b10000000000000000010111100111011; // input=-2.763671875, output=-0.368988769637
			11'd1732: out = 32'b10000000000000000010111011000100; // input=-2.767578125, output=-0.365355362723
			11'd1733: out = 32'b10000000000000000010111001001101; // input=-2.771484375, output=-0.361716380935
			11'd1734: out = 32'b10000000000000000010110111010101; // input=-2.775390625, output=-0.358071879801
			11'd1735: out = 32'b10000000000000000010110101011110; // input=-2.779296875, output=-0.35442191493
			11'd1736: out = 32'b10000000000000000010110011100110; // input=-2.783203125, output=-0.350766542017
			11'd1737: out = 32'b10000000000000000010110001101110; // input=-2.787109375, output=-0.347105816838
			11'd1738: out = 32'b10000000000000000010101111110110; // input=-2.791015625, output=-0.343439795251
			11'd1739: out = 32'b10000000000000000010101101111110; // input=-2.794921875, output=-0.339768533196
			11'd1740: out = 32'b10000000000000000010101100000101; // input=-2.798828125, output=-0.336092086691
			11'd1741: out = 32'b10000000000000000010101010001100; // input=-2.802734375, output=-0.332410511834
			11'd1742: out = 32'b10000000000000000010101000010100; // input=-2.806640625, output=-0.328723864801
			11'd1743: out = 32'b10000000000000000010100110011011; // input=-2.810546875, output=-0.325032201847
			11'd1744: out = 32'b10000000000000000010100100100010; // input=-2.814453125, output=-0.321335579302
			11'd1745: out = 32'b10000000000000000010100010101000; // input=-2.818359375, output=-0.31763405357
			11'd1746: out = 32'b10000000000000000010100000101111; // input=-2.822265625, output=-0.313927681134
			11'd1747: out = 32'b10000000000000000010011110110101; // input=-2.826171875, output=-0.310216518548
			11'd1748: out = 32'b10000000000000000010011100111011; // input=-2.830078125, output=-0.306500622439
			11'd1749: out = 32'b10000000000000000010011011000001; // input=-2.833984375, output=-0.302780049508
			11'd1750: out = 32'b10000000000000000010011001000111; // input=-2.837890625, output=-0.299054856526
			11'd1751: out = 32'b10000000000000000010010111001101; // input=-2.841796875, output=-0.295325100335
			11'd1752: out = 32'b10000000000000000010010101010011; // input=-2.845703125, output=-0.291590837846
			11'd1753: out = 32'b10000000000000000010010011011000; // input=-2.849609375, output=-0.28785212604
			11'd1754: out = 32'b10000000000000000010010001011110; // input=-2.853515625, output=-0.284109021964
			11'd1755: out = 32'b10000000000000000010001111100011; // input=-2.857421875, output=-0.280361582734
			11'd1756: out = 32'b10000000000000000010001101101000; // input=-2.861328125, output=-0.276609865532
			11'd1757: out = 32'b10000000000000000010001011101101; // input=-2.865234375, output=-0.272853927603
			11'd1758: out = 32'b10000000000000000010001001110010; // input=-2.869140625, output=-0.269093826259
			11'd1759: out = 32'b10000000000000000010000111110110; // input=-2.873046875, output=-0.265329618874
			11'd1760: out = 32'b10000000000000000010000101111011; // input=-2.876953125, output=-0.261561362886
			11'd1761: out = 32'b10000000000000000010000011111111; // input=-2.880859375, output=-0.257789115793
			11'd1762: out = 32'b10000000000000000010000010000011; // input=-2.884765625, output=-0.254012935156
			11'd1763: out = 32'b10000000000000000010000000001000; // input=-2.888671875, output=-0.250232878593
			11'd1764: out = 32'b10000000000000000001111110001100; // input=-2.892578125, output=-0.246449003785
			11'd1765: out = 32'b10000000000000000001111100010000; // input=-2.896484375, output=-0.242661368468
			11'd1766: out = 32'b10000000000000000001111010010011; // input=-2.900390625, output=-0.238870030437
			11'd1767: out = 32'b10000000000000000001111000010111; // input=-2.904296875, output=-0.235075047543
			11'd1768: out = 32'b10000000000000000001110110011010; // input=-2.908203125, output=-0.231276477694
			11'd1769: out = 32'b10000000000000000001110100011110; // input=-2.912109375, output=-0.22747437885
			11'd1770: out = 32'b10000000000000000001110010100001; // input=-2.916015625, output=-0.223668809027
			11'd1771: out = 32'b10000000000000000001110000100100; // input=-2.919921875, output=-0.219859826292
			11'd1772: out = 32'b10000000000000000001101110100111; // input=-2.923828125, output=-0.216047488768
			11'd1773: out = 32'b10000000000000000001101100101010; // input=-2.927734375, output=-0.212231854624
			11'd1774: out = 32'b10000000000000000001101010101101; // input=-2.931640625, output=-0.208412982084
			11'd1775: out = 32'b10000000000000000001101000110000; // input=-2.935546875, output=-0.204590929418
			11'd1776: out = 32'b10000000000000000001100110110011; // input=-2.939453125, output=-0.200765754946
			11'd1777: out = 32'b10000000000000000001100100110101; // input=-2.943359375, output=-0.196937517036
			11'd1778: out = 32'b10000000000000000001100010111000; // input=-2.947265625, output=-0.193106274101
			11'd1779: out = 32'b10000000000000000001100000111010; // input=-2.951171875, output=-0.189272084602
			11'd1780: out = 32'b10000000000000000001011110111100; // input=-2.955078125, output=-0.185435007044
			11'd1781: out = 32'b10000000000000000001011100111111; // input=-2.958984375, output=-0.181595099977
			11'd1782: out = 32'b10000000000000000001011011000001; // input=-2.962890625, output=-0.177752421991
			11'd1783: out = 32'b10000000000000000001011001000011; // input=-2.966796875, output=-0.173907031722
			11'd1784: out = 32'b10000000000000000001010111000100; // input=-2.970703125, output=-0.170058987846
			11'd1785: out = 32'b10000000000000000001010101000110; // input=-2.974609375, output=-0.166208349078
			11'd1786: out = 32'b10000000000000000001010011001000; // input=-2.978515625, output=-0.162355174176
			11'd1787: out = 32'b10000000000000000001010001001010; // input=-2.982421875, output=-0.158499521934
			11'd1788: out = 32'b10000000000000000001001111001011; // input=-2.986328125, output=-0.154641451184
			11'd1789: out = 32'b10000000000000000001001101001101; // input=-2.990234375, output=-0.150781020795
			11'd1790: out = 32'b10000000000000000001001011001110; // input=-2.994140625, output=-0.146918289674
			11'd1791: out = 32'b10000000000000000001001001010000; // input=-2.998046875, output=-0.14305331676
			11'd1792: out = 32'b10000000000000000001000111010001; // input=-3.001953125, output=-0.139186161029
			11'd1793: out = 32'b10000000000000000001000101010010; // input=-3.005859375, output=-0.135316881489
			11'd1794: out = 32'b10000000000000000001000011010011; // input=-3.009765625, output=-0.131445537179
			11'd1795: out = 32'b10000000000000000001000001010100; // input=-3.013671875, output=-0.127572187172
			11'd1796: out = 32'b10000000000000000000111111010101; // input=-3.017578125, output=-0.12369689057
			11'd1797: out = 32'b10000000000000000000111101010110; // input=-3.021484375, output=-0.119819706506
			11'd1798: out = 32'b10000000000000000000111011010111; // input=-3.025390625, output=-0.115940694141
			11'd1799: out = 32'b10000000000000000000111001011000; // input=-3.029296875, output=-0.112059912663
			11'd1800: out = 32'b10000000000000000000110111011001; // input=-3.033203125, output=-0.108177421289
			11'd1801: out = 32'b10000000000000000000110101011001; // input=-3.037109375, output=-0.10429327926
			11'd1802: out = 32'b10000000000000000000110011011010; // input=-3.041015625, output=-0.100407545845
			11'd1803: out = 32'b10000000000000000000110001011011; // input=-3.044921875, output=-0.0965202803338
			11'd1804: out = 32'b10000000000000000000101111011011; // input=-3.048828125, output=-0.0926315420419
			11'd1805: out = 32'b10000000000000000000101101011100; // input=-3.052734375, output=-0.0887413903066
			11'd1806: out = 32'b10000000000000000000101011011100; // input=-3.056640625, output=-0.0848498844869
			11'd1807: out = 32'b10000000000000000000101001011101; // input=-3.060546875, output=-0.0809570839624
			11'd1808: out = 32'b10000000000000000000100111011101; // input=-3.064453125, output=-0.0770630481324
			11'd1809: out = 32'b10000000000000000000100101011110; // input=-3.068359375, output=-0.0731678364151
			11'd1810: out = 32'b10000000000000000000100011011110; // input=-3.072265625, output=-0.0692715082466
			11'd1811: out = 32'b10000000000000000000100001011110; // input=-3.076171875, output=-0.0653741230801
			11'd1812: out = 32'b10000000000000000000011111011110; // input=-3.080078125, output=-0.061475740385
			11'd1813: out = 32'b10000000000000000000011101011111; // input=-3.083984375, output=-0.0575764196456
			11'd1814: out = 32'b10000000000000000000011011011111; // input=-3.087890625, output=-0.053676220361
			11'd1815: out = 32'b10000000000000000000011001011111; // input=-3.091796875, output=-0.0497752020432
			11'd1816: out = 32'b10000000000000000000010111011111; // input=-3.095703125, output=-0.0458734242172
			11'd1817: out = 32'b10000000000000000000010101011111; // input=-3.099609375, output=-0.0419709464191
			11'd1818: out = 32'b10000000000000000000010011011111; // input=-3.103515625, output=-0.038067828196
			11'd1819: out = 32'b10000000000000000000010001011111; // input=-3.107421875, output=-0.0341641291047
			11'd1820: out = 32'b10000000000000000000001111100000; // input=-3.111328125, output=-0.0302599087108
			11'd1821: out = 32'b10000000000000000000001101100000; // input=-3.115234375, output=-0.0263552265879
			11'd1822: out = 32'b10000000000000000000001011100000; // input=-3.119140625, output=-0.0224501423167
			11'd1823: out = 32'b10000000000000000000001001100000; // input=-3.123046875, output=-0.018544715484
			11'd1824: out = 32'b10000000000000000000000111100000; // input=-3.126953125, output=-0.0146390056817
			11'd1825: out = 32'b10000000000000000000000101100000; // input=-3.130859375, output=-0.0107330725062
			11'd1826: out = 32'b10000000000000000000000011100000; // input=-3.134765625, output=-0.0068269755572
			11'd1827: out = 32'b10000000000000000000000001100000; // input=-3.138671875, output=-0.00292077443696
			11'd1828: out = 32'b00000000000000000000000000100000; // input=-3.142578125, output=0.000985471250699
			11'd1829: out = 32'b00000000000000000000000010100000; // input=-3.146484375, output=0.00489170190128
			11'd1830: out = 32'b00000000000000000000000100100000; // input=-3.150390625, output=0.00879785791051
			11'd1831: out = 32'b00000000000000000000000110100000; // input=-3.154296875, output=0.0127038796752
			11'd1832: out = 32'b00000000000000000000001000100000; // input=-3.158203125, output=0.0166097075944
			11'd1833: out = 32'b00000000000000000000001010100000; // input=-3.162109375, output=0.0205152820699
			11'd1834: out = 32'b00000000000000000000001100100000; // input=-3.166015625, output=0.0244205435074
			11'd1835: out = 32'b00000000000000000000001110100000; // input=-3.169921875, output=0.0283254323174
			11'd1836: out = 32'b00000000000000000000010000100000; // input=-3.173828125, output=0.0322298889162
			11'd1837: out = 32'b00000000000000000000010010100000; // input=-3.177734375, output=0.0361338537266
			11'd1838: out = 32'b00000000000000000000010100100000; // input=-3.181640625, output=0.0400372671788
			11'd1839: out = 32'b00000000000000000000010110100000; // input=-3.185546875, output=0.0439400697116
			11'd1840: out = 32'b00000000000000000000011000100000; // input=-3.189453125, output=0.0478422017729
			11'd1841: out = 32'b00000000000000000000011010100000; // input=-3.193359375, output=0.0517436038212
			11'd1842: out = 32'b00000000000000000000011100011111; // input=-3.197265625, output=0.0556442163256
			11'd1843: out = 32'b00000000000000000000011110011111; // input=-3.201171875, output=0.0595439797679
			11'd1844: out = 32'b00000000000000000000100000011111; // input=-3.205078125, output=0.0634428346422
			11'd1845: out = 32'b00000000000000000000100010011111; // input=-3.208984375, output=0.0673407214569
			11'd1846: out = 32'b00000000000000000000100100011110; // input=-3.212890625, output=0.0712375807351
			11'd1847: out = 32'b00000000000000000000100110011110; // input=-3.216796875, output=0.0751333530155
			11'd1848: out = 32'b00000000000000000000101000011110; // input=-3.220703125, output=0.0790279788533
			11'd1849: out = 32'b00000000000000000000101010011101; // input=-3.224609375, output=0.0829213988214
			11'd1850: out = 32'b00000000000000000000101100011101; // input=-3.228515625, output=0.086813553511
			11'd1851: out = 32'b00000000000000000000101110011100; // input=-3.232421875, output=0.0907043835325
			11'd1852: out = 32'b00000000000000000000110000011100; // input=-3.236328125, output=0.0945938295168
			11'd1853: out = 32'b00000000000000000000110010011011; // input=-3.240234375, output=0.0984818321156
			11'd1854: out = 32'b00000000000000000000110100011010; // input=-3.244140625, output=0.102368332003
			11'd1855: out = 32'b00000000000000000000110110011010; // input=-3.248046875, output=0.106253269875
			11'd1856: out = 32'b00000000000000000000111000011001; // input=-3.251953125, output=0.110136586453
			11'd1857: out = 32'b00000000000000000000111010011000; // input=-3.255859375, output=0.114018222483
			11'd1858: out = 32'b00000000000000000000111100010111; // input=-3.259765625, output=0.117898118735
			11'd1859: out = 32'b00000000000000000000111110010110; // input=-3.263671875, output=0.121776216006
			11'd1860: out = 32'b00000000000000000001000000010101; // input=-3.267578125, output=0.125652455122
			11'd1861: out = 32'b00000000000000000001000010010100; // input=-3.271484375, output=0.129526776936
			11'd1862: out = 32'b00000000000000000001000100010011; // input=-3.275390625, output=0.133399122331
			11'd1863: out = 32'b00000000000000000001000110010010; // input=-3.279296875, output=0.13726943222
			11'd1864: out = 32'b00000000000000000001001000010001; // input=-3.283203125, output=0.141137647546
			11'd1865: out = 32'b00000000000000000001001010001111; // input=-3.287109375, output=0.145003709285
			11'd1866: out = 32'b00000000000000000001001100001110; // input=-3.291015625, output=0.148867558446
			11'd1867: out = 32'b00000000000000000001001110001101; // input=-3.294921875, output=0.152729136071
			11'd1868: out = 32'b00000000000000000001010000001011; // input=-3.298828125, output=0.156588383237
			11'd1869: out = 32'b00000000000000000001010010001001; // input=-3.302734375, output=0.160445241058
			11'd1870: out = 32'b00000000000000000001010100001000; // input=-3.306640625, output=0.164299650681
			11'd1871: out = 32'b00000000000000000001010110000110; // input=-3.310546875, output=0.168151553294
			11'd1872: out = 32'b00000000000000000001011000000100; // input=-3.314453125, output=0.172000890121
			11'd1873: out = 32'b00000000000000000001011010000010; // input=-3.318359375, output=0.175847602426
			11'd1874: out = 32'b00000000000000000001011100000000; // input=-3.322265625, output=0.179691631513
			11'd1875: out = 32'b00000000000000000001011101111110; // input=-3.326171875, output=0.183532918727
			11'd1876: out = 32'b00000000000000000001011111111100; // input=-3.330078125, output=0.187371405454
			11'd1877: out = 32'b00000000000000000001100001111001; // input=-3.333984375, output=0.191207033124
			11'd1878: out = 32'b00000000000000000001100011110111; // input=-3.337890625, output=0.19503974321
			11'd1879: out = 32'b00000000000000000001100101110101; // input=-3.341796875, output=0.198869477229
			11'd1880: out = 32'b00000000000000000001100111110010; // input=-3.345703125, output=0.202696176745
			11'd1881: out = 32'b00000000000000000001101001101111; // input=-3.349609375, output=0.206519783367
			11'd1882: out = 32'b00000000000000000001101011101100; // input=-3.353515625, output=0.210340238751
			11'd1883: out = 32'b00000000000000000001101101101010; // input=-3.357421875, output=0.214157484602
			11'd1884: out = 32'b00000000000000000001101111100110; // input=-3.361328125, output=0.217971462672
			11'd1885: out = 32'b00000000000000000001110001100011; // input=-3.365234375, output=0.221782114767
			11'd1886: out = 32'b00000000000000000001110011100000; // input=-3.369140625, output=0.225589382739
			11'd1887: out = 32'b00000000000000000001110101011101; // input=-3.373046875, output=0.229393208495
			11'd1888: out = 32'b00000000000000000001110111011001; // input=-3.376953125, output=0.233193533993
			11'd1889: out = 32'b00000000000000000001111001010110; // input=-3.380859375, output=0.236990301245
			11'd1890: out = 32'b00000000000000000001111011010010; // input=-3.384765625, output=0.240783452315
			11'd1891: out = 32'b00000000000000000001111101001110; // input=-3.388671875, output=0.244572929327
			11'd1892: out = 32'b00000000000000000001111111001010; // input=-3.392578125, output=0.248358674457
			11'd1893: out = 32'b00000000000000000010000001000110; // input=-3.396484375, output=0.252140629939
			11'd1894: out = 32'b00000000000000000010000011000010; // input=-3.400390625, output=0.255918738065
			11'd1895: out = 32'b00000000000000000010000100111110; // input=-3.404296875, output=0.259692941186
			11'd1896: out = 32'b00000000000000000010000110111001; // input=-3.408203125, output=0.263463181712
			11'd1897: out = 32'b00000000000000000010001000110101; // input=-3.412109375, output=0.267229402115
			11'd1898: out = 32'b00000000000000000010001010110000; // input=-3.416015625, output=0.270991544925
			11'd1899: out = 32'b00000000000000000010001100101011; // input=-3.419921875, output=0.274749552738
			11'd1900: out = 32'b00000000000000000010001110100110; // input=-3.423828125, output=0.27850336821
			11'd1901: out = 32'b00000000000000000010010000100001; // input=-3.427734375, output=0.282252934064
			11'd1902: out = 32'b00000000000000000010010010011100; // input=-3.431640625, output=0.285998193086
			11'd1903: out = 32'b00000000000000000010010100010110; // input=-3.435546875, output=0.289739088127
			11'd1904: out = 32'b00000000000000000010010110010001; // input=-3.439453125, output=0.293475562106
			11'd1905: out = 32'b00000000000000000010011000001011; // input=-3.443359375, output=0.297207558008
			11'd1906: out = 32'b00000000000000000010011010000101; // input=-3.447265625, output=0.30093501889
			11'd1907: out = 32'b00000000000000000010011011111111; // input=-3.451171875, output=0.304657887873
			11'd1908: out = 32'b00000000000000000010011101111001; // input=-3.455078125, output=0.308376108151
			11'd1909: out = 32'b00000000000000000010011111110011; // input=-3.458984375, output=0.31208962299
			11'd1910: out = 32'b00000000000000000010100001101100; // input=-3.462890625, output=0.315798375725
			11'd1911: out = 32'b00000000000000000010100011100101; // input=-3.466796875, output=0.319502309765
			11'd1912: out = 32'b00000000000000000010100101011111; // input=-3.470703125, output=0.323201368593
			11'd1913: out = 32'b00000000000000000010100111011000; // input=-3.474609375, output=0.326895495766
			11'd1914: out = 32'b00000000000000000010101001010001; // input=-3.478515625, output=0.330584634915
			11'd1915: out = 32'b00000000000000000010101011001001; // input=-3.482421875, output=0.33426872975
			11'd1916: out = 32'b00000000000000000010101101000010; // input=-3.486328125, output=0.337947724056
			11'd1917: out = 32'b00000000000000000010101110111010; // input=-3.490234375, output=0.341621561694
			11'd1918: out = 32'b00000000000000000010110000110010; // input=-3.494140625, output=0.345290186609
			11'd1919: out = 32'b00000000000000000010110010101011; // input=-3.498046875, output=0.348953542819
			11'd1920: out = 32'b00000000000000000010110100100010; // input=-3.501953125, output=0.352611574428
			11'd1921: out = 32'b00000000000000000010110110011010; // input=-3.505859375, output=0.356264225619
			11'd1922: out = 32'b00000000000000000010111000010010; // input=-3.509765625, output=0.359911440655
			11'd1923: out = 32'b00000000000000000010111010001001; // input=-3.513671875, output=0.363553163886
			11'd1924: out = 32'b00000000000000000010111100000000; // input=-3.517578125, output=0.367189339743
			11'd1925: out = 32'b00000000000000000010111101110111; // input=-3.521484375, output=0.370819912742
			11'd1926: out = 32'b00000000000000000010111111101110; // input=-3.525390625, output=0.374444827485
			11'd1927: out = 32'b00000000000000000011000001100100; // input=-3.529296875, output=0.378064028661
			11'd1928: out = 32'b00000000000000000011000011011011; // input=-3.533203125, output=0.381677461046
			11'd1929: out = 32'b00000000000000000011000101010001; // input=-3.537109375, output=0.385285069501
			11'd1930: out = 32'b00000000000000000011000111000111; // input=-3.541015625, output=0.388886798981
			11'd1931: out = 32'b00000000000000000011001000111101; // input=-3.544921875, output=0.392482594526
			11'd1932: out = 32'b00000000000000000011001010110011; // input=-3.548828125, output=0.39607240127
			11'd1933: out = 32'b00000000000000000011001100101000; // input=-3.552734375, output=0.399656164437
			11'd1934: out = 32'b00000000000000000011001110011101; // input=-3.556640625, output=0.403233829342
			11'd1935: out = 32'b00000000000000000011010000010010; // input=-3.560546875, output=0.406805341395
			11'd1936: out = 32'b00000000000000000011010010000111; // input=-3.564453125, output=0.410370646099
			11'd1937: out = 32'b00000000000000000011010011111100; // input=-3.568359375, output=0.413929689052
			11'd1938: out = 32'b00000000000000000011010101110000; // input=-3.572265625, output=0.417482415947
			11'd1939: out = 32'b00000000000000000011010111100100; // input=-3.576171875, output=0.421028772574
			11'd1940: out = 32'b00000000000000000011011001011000; // input=-3.580078125, output=0.42456870482
			11'd1941: out = 32'b00000000000000000011011011001100; // input=-3.583984375, output=0.42810215867
			11'd1942: out = 32'b00000000000000000011011101000000; // input=-3.587890625, output=0.431629080208
			11'd1943: out = 32'b00000000000000000011011110110011; // input=-3.591796875, output=0.435149415617
			11'd1944: out = 32'b00000000000000000011100000100110; // input=-3.595703125, output=0.438663111181
			11'd1945: out = 32'b00000000000000000011100010011001; // input=-3.599609375, output=0.442170113286
			11'd1946: out = 32'b00000000000000000011100100001100; // input=-3.603515625, output=0.445670368419
			11'd1947: out = 32'b00000000000000000011100101111110; // input=-3.607421875, output=0.44916382317
			11'd1948: out = 32'b00000000000000000011100111110000; // input=-3.611328125, output=0.452650424234
			11'd1949: out = 32'b00000000000000000011101001100010; // input=-3.615234375, output=0.45613011841
			11'd1950: out = 32'b00000000000000000011101011010100; // input=-3.619140625, output=0.459602852601
			11'd1951: out = 32'b00000000000000000011101101000110; // input=-3.623046875, output=0.463068573818
			11'd1952: out = 32'b00000000000000000011101110110111; // input=-3.626953125, output=0.466527229179
			11'd1953: out = 32'b00000000000000000011110000101000; // input=-3.630859375, output=0.469978765908
			11'd1954: out = 32'b00000000000000000011110010011001; // input=-3.634765625, output=0.473423131339
			11'd1955: out = 32'b00000000000000000011110100001010; // input=-3.638671875, output=0.476860272915
			11'd1956: out = 32'b00000000000000000011110101111010; // input=-3.642578125, output=0.480290138191
			11'd1957: out = 32'b00000000000000000011110111101010; // input=-3.646484375, output=0.48371267483
			11'd1958: out = 32'b00000000000000000011111001011010; // input=-3.650390625, output=0.487127830609
			11'd1959: out = 32'b00000000000000000011111011001010; // input=-3.654296875, output=0.490535553416
			11'd1960: out = 32'b00000000000000000011111100111001; // input=-3.658203125, output=0.493935791254
			11'd1961: out = 32'b00000000000000000011111110101000; // input=-3.662109375, output=0.49732849224
			11'd1962: out = 32'b00000000000000000100000000010111; // input=-3.666015625, output=0.500713604605
			11'd1963: out = 32'b00000000000000000100000010000110; // input=-3.669921875, output=0.504091076697
			11'd1964: out = 32'b00000000000000000100000011110100; // input=-3.673828125, output=0.507460856978
			11'd1965: out = 32'b00000000000000000100000101100011; // input=-3.677734375, output=0.510822894032
			11'd1966: out = 32'b00000000000000000100000111010001; // input=-3.681640625, output=0.514177136557
			11'd1967: out = 32'b00000000000000000100001000111110; // input=-3.685546875, output=0.517523533371
			11'd1968: out = 32'b00000000000000000100001010101100; // input=-3.689453125, output=0.520862033412
			11'd1969: out = 32'b00000000000000000100001100011001; // input=-3.693359375, output=0.52419258574
			11'd1970: out = 32'b00000000000000000100001110000110; // input=-3.697265625, output=0.527515139534
			11'd1971: out = 32'b00000000000000000100001111110010; // input=-3.701171875, output=0.530829644096
			11'd1972: out = 32'b00000000000000000100010001011111; // input=-3.705078125, output=0.534136048851
			11'd1973: out = 32'b00000000000000000100010011001011; // input=-3.708984375, output=0.537434303347
			11'd1974: out = 32'b00000000000000000100010100110110; // input=-3.712890625, output=0.540724357256
			11'd1975: out = 32'b00000000000000000100010110100010; // input=-3.716796875, output=0.544006160377
			11'd1976: out = 32'b00000000000000000100011000001101; // input=-3.720703125, output=0.547279662634
			11'd1977: out = 32'b00000000000000000100011001111000; // input=-3.724609375, output=0.550544814076
			11'd1978: out = 32'b00000000000000000100011011100011; // input=-3.728515625, output=0.553801564881
			11'd1979: out = 32'b00000000000000000100011101001101; // input=-3.732421875, output=0.557049865356
			11'd1980: out = 32'b00000000000000000100011110111000; // input=-3.736328125, output=0.560289665936
			11'd1981: out = 32'b00000000000000000100100000100001; // input=-3.740234375, output=0.563520917184
			11'd1982: out = 32'b00000000000000000100100010001011; // input=-3.744140625, output=0.566743569797
			11'd1983: out = 32'b00000000000000000100100011110100; // input=-3.748046875, output=0.5699575746
			11'd1984: out = 32'b00000000000000000100100101011101; // input=-3.751953125, output=0.573162882552
			11'd1985: out = 32'b00000000000000000100100111000110; // input=-3.755859375, output=0.576359444743
			11'd1986: out = 32'b00000000000000000100101000101111; // input=-3.759765625, output=0.579547212398
			11'd1987: out = 32'b00000000000000000100101010010111; // input=-3.763671875, output=0.582726136876
			11'd1988: out = 32'b00000000000000000100101011111111; // input=-3.767578125, output=0.58589616967
			11'd1989: out = 32'b00000000000000000100101101100110; // input=-3.771484375, output=0.58905726241
			11'd1990: out = 32'b00000000000000000100101111001110; // input=-3.775390625, output=0.59220936686
			11'd1991: out = 32'b00000000000000000100110000110101; // input=-3.779296875, output=0.595352434924
			11'd1992: out = 32'b00000000000000000100110010011011; // input=-3.783203125, output=0.598486418642
			11'd1993: out = 32'b00000000000000000100110100000010; // input=-3.787109375, output=0.601611270194
			11'd1994: out = 32'b00000000000000000100110101101000; // input=-3.791015625, output=0.604726941898
			11'd1995: out = 32'b00000000000000000100110111001101; // input=-3.794921875, output=0.607833386213
			11'd1996: out = 32'b00000000000000000100111000110011; // input=-3.798828125, output=0.610930555738
			11'd1997: out = 32'b00000000000000000100111010011000; // input=-3.802734375, output=0.614018403215
			11'd1998: out = 32'b00000000000000000100111011111101; // input=-3.806640625, output=0.617096881526
			11'd1999: out = 32'b00000000000000000100111101100010; // input=-3.810546875, output=0.620165943698
			11'd2000: out = 32'b00000000000000000100111111000110; // input=-3.814453125, output=0.623225542901
			11'd2001: out = 32'b00000000000000000101000000101010; // input=-3.818359375, output=0.626275632449
			11'd2002: out = 32'b00000000000000000101000010001101; // input=-3.822265625, output=0.629316165801
			11'd2003: out = 32'b00000000000000000101000011110001; // input=-3.826171875, output=0.632347096563
			11'd2004: out = 32'b00000000000000000101000101010100; // input=-3.830078125, output=0.635368378486
			11'd2005: out = 32'b00000000000000000101000110110110; // input=-3.833984375, output=0.638379965469
			11'd2006: out = 32'b00000000000000000101001000011001; // input=-3.837890625, output=0.64138181156
			11'd2007: out = 32'b00000000000000000101001001111011; // input=-3.841796875, output=0.644373870953
			11'd2008: out = 32'b00000000000000000101001011011101; // input=-3.845703125, output=0.647356097993
			11'd2009: out = 32'b00000000000000000101001100111110; // input=-3.849609375, output=0.650328447176
			11'd2010: out = 32'b00000000000000000101001110011111; // input=-3.853515625, output=0.653290873148
			11'd2011: out = 32'b00000000000000000101010000000000; // input=-3.857421875, output=0.656243330704
			11'd2012: out = 32'b00000000000000000101010001100000; // input=-3.861328125, output=0.659185774794
			11'd2013: out = 32'b00000000000000000101010011000000; // input=-3.865234375, output=0.662118160521
			11'd2014: out = 32'b00000000000000000101010100100000; // input=-3.869140625, output=0.665040443139
			11'd2015: out = 32'b00000000000000000101010101111111; // input=-3.873046875, output=0.667952578058
			11'd2016: out = 32'b00000000000000000101010111011111; // input=-3.876953125, output=0.670854520842
			11'd2017: out = 32'b00000000000000000101011000111101; // input=-3.880859375, output=0.673746227212
			11'd2018: out = 32'b00000000000000000101011010011100; // input=-3.884765625, output=0.676627653043
			11'd2019: out = 32'b00000000000000000101011011111010; // input=-3.888671875, output=0.679498754369
			11'd2020: out = 32'b00000000000000000101011101011000; // input=-3.892578125, output=0.68235948738
			11'd2021: out = 32'b00000000000000000101011110110101; // input=-3.896484375, output=0.685209808425
			11'd2022: out = 32'b00000000000000000101100000010010; // input=-3.900390625, output=0.688049674011
			11'd2023: out = 32'b00000000000000000101100001101111; // input=-3.904296875, output=0.690879040805
			11'd2024: out = 32'b00000000000000000101100011001011; // input=-3.908203125, output=0.693697865636
			11'd2025: out = 32'b00000000000000000101100100100111; // input=-3.912109375, output=0.69650610549
			11'd2026: out = 32'b00000000000000000101100110000011; // input=-3.916015625, output=0.699303717518
			11'd2027: out = 32'b00000000000000000101100111011110; // input=-3.919921875, output=0.702090659032
			11'd2028: out = 32'b00000000000000000101101000111001; // input=-3.923828125, output=0.704866887506
			11'd2029: out = 32'b00000000000000000101101010010100; // input=-3.927734375, output=0.707632360579
			11'd2030: out = 32'b00000000000000000101101011101110; // input=-3.931640625, output=0.710387036053
			11'd2031: out = 32'b00000000000000000101101101001000; // input=-3.935546875, output=0.713130871894
			11'd2032: out = 32'b00000000000000000101101110100001; // input=-3.939453125, output=0.715863826236
			11'd2033: out = 32'b00000000000000000101101111111011; // input=-3.943359375, output=0.718585857376
			11'd2034: out = 32'b00000000000000000101110001010011; // input=-3.947265625, output=0.72129692378
			11'd2035: out = 32'b00000000000000000101110010101100; // input=-3.951171875, output=0.723996984081
			11'd2036: out = 32'b00000000000000000101110100000100; // input=-3.955078125, output=0.726685997079
			11'd2037: out = 32'b00000000000000000101110101011100; // input=-3.958984375, output=0.729363921742
			11'd2038: out = 32'b00000000000000000101110110110011; // input=-3.962890625, output=0.732030717209
			11'd2039: out = 32'b00000000000000000101111000001010; // input=-3.966796875, output=0.734686342788
			11'd2040: out = 32'b00000000000000000101111001100001; // input=-3.970703125, output=0.737330757958
			11'd2041: out = 32'b00000000000000000101111010110111; // input=-3.974609375, output=0.739963922367
			11'd2042: out = 32'b00000000000000000101111100001101; // input=-3.978515625, output=0.742585795837
			11'd2043: out = 32'b00000000000000000101111101100011; // input=-3.982421875, output=0.745196338362
			11'd2044: out = 32'b00000000000000000101111110111000; // input=-3.986328125, output=0.747795510107
			11'd2045: out = 32'b00000000000000000110000000001101; // input=-3.990234375, output=0.750383271413
			11'd2046: out = 32'b00000000000000000110000001100001; // input=-3.994140625, output=0.752959582793
			11'd2047: out = 32'b00000000000000000110000010110101; // input=-3.998046875, output=0.755524404937
		endcase
	end
	converter U0 (a, index);

endmodule

module converter(a, index);
	input  [31:0] a;
	output [10:0] index;

	assign index[10]	= a[31];
	assign index[9:8]	= a[16:15];
	assign index[7:0]	= a[14:7];
endmodule
