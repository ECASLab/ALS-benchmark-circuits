`timescale 1ns / 1ps

module RForest(
	A1,
	A2,
	A3,
	A4,
	A5,
	A6,
	A7,
	A8,
	A9,
	A91,
	A92,
	A93,
	A94,
	A95,
	A96,
	A97,
	A98,
	A99,
	A991,
	A992,
	A993,
	A994,
	A995,
	A996,
	A997,
	A998,
	A999,
	A9991,
	A9992,
	A9993,
	A9994,
	A9995,
	A9996,
	A9997,
	A9998,
	A9999,
	A99991,
	A99992,
	A99993,
	A99994,
	A99995,
	A99996,
	A99997,
	A99998,
	A99999,
	A999991,
	A999992,
	A999993,
	A999994,
	A999995,
	A999996,
	A999997,
	decision
);


	input [9:0] A1;
	input [9:0] A2;
	input [9:0] A3;
	input [9:0] A4;
	input [9:0] A5;
	input [9:0] A6;
	input [9:0] A7;
	input [9:0] A8;
	input [9:0] A9;
	input [9:0] A91;
	input [9:0] A92;
	input [9:0] A93;
	input [9:0] A94;
	input [9:0] A95;
	input [9:0] A96;
	input [9:0] A97;
	input [9:0] A98;
	input [9:0] A99;
	input [9:0] A991;
	input [9:0] A992;
	input [9:0] A993;
	input [9:0] A994;
	input [9:0] A995;
	input [9:0] A996;
	input [9:0] A997;
	input [9:0] A998;
	input [9:0] A999;
	input [9:0] A9991;
	input [9:0] A9992;
	input [9:0] A9993;
	input [9:0] A9994;
	input [9:0] A9995;
	input [9:0] A9996;
	input [9:0] A9997;
	input [9:0] A9998;
	input [9:0] A9999;
	input [9:0] A99991;
	input [9:0] A99992;
	input [9:0] A99993;
	input [9:0] A99994;
	input [9:0] A99995;
	input [9:0] A99996;
	input [9:0] A99997;
	input [9:0] A99998;
	input [9:0] A99999;
	input [9:0] A999991;
	input [9:0] A999992;
	input [9:0] A999993;
	input [9:0] A999994;
	input [9:0] A999995;
	input [9:0] A999996;
	input [9:0] A999997;
	output [4:0] decision;

	wire [9:0] reg_A1;
	wire [9:0] reg_A2;
	wire [9:0] reg_A3;
	wire [9:0] reg_A4;
	wire [9:0] reg_A5;
	wire [9:0] reg_A6;
	wire [9:0] reg_A7;
	wire [9:0] reg_A8;
	wire [9:0] reg_A9;
	wire [9:0] reg_A91;
	wire [9:0] reg_A92;
	wire [9:0] reg_A93;
	wire [9:0] reg_A94;
	wire [9:0] reg_A95;
	wire [9:0] reg_A96;
	wire [9:0] reg_A97;
	wire [9:0] reg_A98;
	wire [9:0] reg_A99;
	wire [9:0] reg_A991;
	wire [9:0] reg_A992;
	wire [9:0] reg_A993;
	wire [9:0] reg_A994;
	wire [9:0] reg_A995;
	wire [9:0] reg_A996;
	wire [9:0] reg_A997;
	wire [9:0] reg_A998;
	wire [9:0] reg_A999;
	wire [9:0] reg_A9991;
	wire [9:0] reg_A9992;
	wire [9:0] reg_A9993;
	wire [9:0] reg_A9994;
	wire [9:0] reg_A9995;
	wire [9:0] reg_A9996;
	wire [9:0] reg_A9997;
	wire [9:0] reg_A9998;
	wire [9:0] reg_A9999;
	wire [9:0] reg_A99991;
	wire [9:0] reg_A99992;
	wire [9:0] reg_A99993;
	wire [9:0] reg_A99994;
	wire [9:0] reg_A99995;
	wire [9:0] reg_A99996;
	wire [9:0] reg_A99997;
	wire [9:0] reg_A99998;
	wire [9:0] reg_A99999;
	wire [9:0] reg_A999991;
	wire [9:0] reg_A999992;
	wire [9:0] reg_A999993;
	wire [9:0] reg_A999994;
	wire [9:0] reg_A999995;
	wire [9:0] reg_A999996;
	wire [9:0] reg_A999997;
	wire [4:0] reg_decision;

wire [0:0] comp_A1_649;
wire [0:0] comp_A2_29;
wire [0:0] comp_A3_322;
wire [0:0] comp_A4_504;
wire [0:0] comp_A5_495;
wire [0:0] comp_A6_624;
wire [0:0] comp_A7_593;
wire [0:0] comp_A1_220;
wire [0:0] comp_A4_472;
wire [0:0] comp_A8_701;
wire [0:0] comp_A9_178;
wire [0:0] comp_A91_362;
wire [0:0] comp_A92_263;
wire [0:0] comp_A93_529;
wire [0:0] comp_A94_40;
wire [0:0] comp_A7_795;
wire [0:0] comp_A95_118;
wire [0:0] comp_A3_541;
wire [0:0] comp_A8_90;
wire [0:0] comp_A96_11;
wire [0:0] comp_A97_193;
wire [0:0] comp_A98_202;
wire [0:0] comp_A99_14;
wire [0:0] comp_A2_830;
wire [0:0] comp_A991_288;
wire [0:0] comp_A992_452;
wire [0:0] comp_A95_373;
wire [0:0] comp_A8_777;
wire [0:0] comp_A93_537;
wire [0:0] comp_A99_11;
wire [0:0] comp_A95_383;
wire [0:0] comp_A993_454;
wire [0:0] comp_A992_774;
wire [0:0] comp_A994_302;
wire [0:0] comp_A995_87;
wire [0:0] comp_A98_143;
wire [0:0] comp_A996_348;
wire [0:0] comp_A997_750;
wire [0:0] comp_A1_884;
wire [0:0] comp_A997_360;
wire [0:0] comp_A998_765;
wire [0:0] comp_A8_726;
wire [0:0] comp_A999_643;
wire [0:0] comp_A3_526;
wire [0:0] comp_A7_455;
wire [0:0] comp_A9991_920;
wire [0:0] comp_A3_300;
wire [0:0] comp_A92_262;
wire [0:0] comp_A9992_183;
wire [0:0] comp_A991_737;
wire [0:0] comp_A97_140;
wire [0:0] comp_A9991_923;
wire [0:0] comp_A96_873;
wire [0:0] comp_A9993_513;
wire [0:0] comp_A4_515;
wire [0:0] comp_A9994_577;
wire [0:0] comp_A94_46;
wire [0:0] comp_A7_341;
wire [0:0] comp_A3_687;
wire [0:0] comp_A9995_483;
wire [0:0] comp_A9996_660;
wire [0:0] comp_A9997_526;
wire [0:0] comp_A9991_943;
wire [0:0] comp_A7_561;
wire [0:0] comp_A993_276;
wire [0:0] comp_A9998_478;
wire [0:0] comp_A92_975;
wire [0:0] comp_A1_727;
wire [0:0] comp_A7_583;
wire [0:0] comp_A995_79;
wire [0:0] comp_A97_173;
wire [0:0] comp_A993_665;
wire [0:0] comp_A9999_801;
wire [0:0] comp_A3_536;
wire [0:0] comp_A999_620;
wire [0:0] comp_A994_700;
wire [0:0] comp_A99991_242;
wire [0:0] comp_A994_712;
wire [0:0] comp_A99992_806;
wire [0:0] comp_A9997_570;
wire [0:0] comp_A99993_119;
wire [0:0] comp_A6_670;
wire [0:0] comp_A994_338;
wire [0:0] comp_A6_635;
wire [0:0] comp_A9994_627;
wire [0:0] comp_A1_881;
wire [0:0] comp_A4_490;
wire [0:0] comp_A92_264;
wire [0:0] comp_A2_839;
wire [0:0] comp_A991_760;
wire [0:0] comp_A993_680;
wire [0:0] comp_A99994_810;
wire [0:0] comp_A98_974;
wire [0:0] comp_A4_350;
wire [0:0] comp_A1_738;
wire [0:0] comp_A997_319;
wire [0:0] comp_A7_411;
wire [0:0] comp_A4_400;
wire [0:0] comp_A9992_93;
wire [0:0] comp_A99994_781;
wire [0:0] comp_A93_726;
wire [0:0] comp_A9998_769;
wire [0:0] comp_A7_415;
wire [0:0] comp_A9991_972;
wire [0:0] comp_A993_608;
wire [0:0] comp_A3_284;
wire [0:0] comp_A9995_876;
wire [0:0] comp_A9_859;
wire [0:0] comp_A9992_129;
wire [0:0] comp_A3_102;
wire [0:0] comp_A3_79;
wire [0:0] comp_A9993_585;
wire [0:0] comp_A3_124;
wire [0:0] comp_A91_239;
wire [0:0] comp_A93_116;
wire [0:0] comp_A9_811;
wire [0:0] comp_A3_757;
wire [0:0] comp_A99991_336;
wire [0:0] comp_A98_66;
wire [0:0] comp_A99995_631;
wire [0:0] comp_A999_732;
wire [0:0] comp_A9996_244;
wire [0:0] comp_A995_167;
wire [0:0] comp_A98_171;
wire [0:0] comp_A3_981;
wire [0:0] comp_A9_827;
wire [0:0] comp_A9992_357;
wire [0:0] comp_A4_739;
wire [0:0] comp_A2_876;
wire [0:0] comp_A99996_412;
wire [0:0] comp_A9996_202;
wire [0:0] comp_A9993_525;
wire [0:0] comp_A7_666;
wire [0:0] comp_A92_519;
wire [0:0] comp_A99994_745;
wire [0:0] comp_A998_448;
wire [0:0] comp_A9997_490;
wire [0:0] comp_A9996_448;
wire [0:0] comp_A997_332;
wire [0:0] comp_A4_495;
wire [0:0] comp_A94_29;
wire [0:0] comp_A7_919;
wire [0:0] comp_A99997_247;
wire [0:0] comp_A993_764;
wire [0:0] comp_A9991_914;
wire [0:0] comp_A96_609;
wire [0:0] comp_A9999_832;
wire [0:0] comp_A99998_189;
wire [0:0] comp_A996_296;
wire [0:0] comp_A99999_409;
wire [0:0] comp_A99994_713;
wire [0:0] comp_A993_839;
wire [0:0] comp_A99997_833;
wire [0:0] comp_A5_327;
wire [0:0] comp_A2_894;
wire [0:0] comp_A3_587;
wire [0:0] comp_A93_629;
wire [0:0] comp_A999991_302;
wire [0:0] comp_A99997_824;
wire [0:0] comp_A9_155;
wire [0:0] comp_A5_170;
wire [0:0] comp_A97_991;
wire [0:0] comp_A995_114;
wire [0:0] comp_A5_586;
wire [0:0] comp_A98_162;
wire [0:0] comp_A991_728;
wire [0:0] comp_A9996_782;
wire [0:0] comp_A99992_505;
wire [0:0] comp_A9995_733;
wire [0:0] comp_A9991_1016;
wire [0:0] comp_A9_152;
wire [0:0] comp_A5_126;
wire [0:0] comp_A999992_426;
wire [0:0] comp_A9_784;
wire [0:0] comp_A999992_487;
wire [0:0] comp_A92_504;
wire [0:0] comp_A9994_769;
wire [0:0] comp_A95_435;
wire [0:0] comp_A999992_569;
wire [0:0] comp_A1_652;
wire [0:0] comp_A991_268;
wire [0:0] comp_A99997_799;
wire [0:0] comp_A992_599;
wire [0:0] comp_A99991_539;
wire [0:0] comp_A98_147;
wire [0:0] comp_A7_591;
wire [0:0] comp_A997_589;
wire [0:0] comp_A97_124;
wire [0:0] comp_A996_225;
wire [0:0] comp_A97_121;
wire [0:0] comp_A99995_671;
wire [0:0] comp_A9998_723;
wire [0:0] comp_A999993_9;
wire [0:0] comp_A996_92;
wire [0:0] comp_A996_222;
wire [0:0] comp_A9999_756;
wire [0:0] comp_A95_203;
wire [0:0] comp_A997_838;
wire [0:0] comp_A5_478;
wire [0:0] comp_A99997_254;
wire [0:0] comp_A99991_618;
wire [0:0] comp_A91_963;
wire [0:0] comp_A9994_288;
wire [0:0] comp_A9991_935;
wire [0:0] comp_A99997_931;
wire [0:0] comp_A98_151;
wire [0:0] comp_A4_486;
wire [0:0] comp_A3_232;
wire [0:0] comp_A9995_839;
wire [0:0] comp_A7_592;
wire [0:0] comp_A3_286;
wire [0:0] comp_A99999_486;
wire [0:0] comp_A9991_932;
wire [0:0] comp_A996_372;
wire [0:0] comp_A9_156;
wire [0:0] comp_A7_804;
wire [0:0] comp_A6_255;
wire [0:0] comp_A99991_344;
wire [0:0] comp_A8_757;
wire [0:0] comp_A993_555;
wire [0:0] comp_A999994_442;
wire [0:0] comp_A99992_671;
wire [0:0] comp_A991_479;
wire [0:0] comp_A97_610;
wire [0:0] comp_A999991_570;
wire [0:0] comp_A9_816;
wire [0:0] comp_A3_80;
wire [0:0] comp_A8_822;
wire [0:0] comp_A998_424;
wire [0:0] comp_A999993_8;
wire [0:0] comp_A9992_421;
wire [0:0] comp_A99999_549;
wire [0:0] comp_A9993_307;
wire [0:0] comp_A9996_562;
wire [0:0] comp_A996_271;
wire [0:0] comp_A992_400;
wire [0:0] comp_A94_31;
wire [0:0] comp_A99_8;
wire [0:0] comp_A3_54;
wire [0:0] comp_A2_872;
wire [0:0] comp_A92_972;
wire [0:0] comp_A3_272;
wire [0:0] comp_A999995_1015;
wire [0:0] comp_A7_605;
wire [0:0] comp_A9993_295;
wire [0:0] comp_A991_531;
wire [0:0] comp_A993_317;
wire [0:0] comp_A991_869;
wire [0:0] comp_A94_50;
wire [0:0] comp_A99994_178;
wire [0:0] comp_A8_786;
wire [0:0] comp_A3_407;
wire [0:0] comp_A6_722;
wire [0:0] comp_A99999_735;
wire [0:0] comp_A92_259;
wire [0:0] comp_A999996_390;
wire [0:0] comp_A2_901;
wire [0:0] comp_A992_675;
wire [0:0] comp_A9_821;
wire [0:0] comp_A92_503;
wire [0:0] comp_A8_536;
wire [0:0] comp_A2_124;
wire [0:0] comp_A92_250;
wire [0:0] comp_A95_497;
wire [0:0] comp_A6_406;
wire [0:0] comp_A9991_948;
wire [0:0] comp_A9999_819;
wire [0:0] comp_A3_535;
wire [0:0] comp_A998_805;
wire [0:0] comp_A92_995;
wire [0:0] comp_A9996_600;
wire [0:0] comp_A6_606;
wire [0:0] comp_A996_353;
wire [0:0] comp_A99994_600;
wire [0:0] comp_A99991_286;
wire [0:0] comp_A996_340;
wire [0:0] comp_A998_414;
wire [0:0] comp_A996_331;
wire [0:0] comp_A994_640;
wire [0:0] comp_A999_714;
wire [0:0] comp_A3_233;
wire [0:0] comp_A9_805;
wire [0:0] comp_A8_540;
wire [0:0] comp_A99996_575;
wire [0:0] comp_A993_982;
wire [0:0] comp_A9993_530;
wire [0:0] comp_A994_475;
wire [0:0] comp_A996_332;
wire [0:0] comp_A4_484;
wire [0:0] comp_A98_325;
wire [0:0] comp_A993_659;
wire [0:0] comp_A2_602;
wire [0:0] comp_A92_505;
wire [0:0] comp_A99999_58;
wire [0:0] comp_A9992_123;
wire [0:0] comp_A999992_527;
wire [0:0] comp_A9996_758;
wire [0:0] comp_A997_428;
wire [0:0] comp_A3_515;
wire [0:0] comp_A992_389;
wire [0:0] comp_A93_513;
wire [0:0] comp_A99999_558;
wire [0:0] comp_A9992_429;
wire [0:0] comp_A993_440;
wire [0:0] comp_A99996_766;
wire [0:0] comp_A999991_485;
wire [0:0] comp_A9991_1009;
wire [0:0] comp_A99999_594;
wire [0:0] comp_A993_492;
wire [0:0] comp_A96_754;
wire [0:0] comp_A993_321;
wire [0:0] comp_A999_712;
wire [0:0] comp_A997_421;
wire [0:0] comp_A9999_805;
wire [0:0] comp_A995_343;
wire [0:0] comp_A9996_570;
wire [0:0] comp_A5_653;
wire [0:0] comp_A4_445;
wire [0:0] comp_A99995_511;
wire [0:0] comp_A99991_185;
wire [0:0] comp_A99999_517;
wire [0:0] comp_A8_334;
wire [0:0] comp_A9996_737;
wire [0:0] comp_A9_845;
wire [0:0] comp_A997_339;
wire [0:0] comp_A997_243;
wire [0:0] comp_A993_683;
wire [0:0] comp_A994_543;
wire [0:0] comp_A99_13;
wire [0:0] comp_A2_22;
wire [0:0] comp_A96_818;
wire [0:0] comp_A3_350;
wire [0:0] comp_A992_528;
wire [0:0] comp_A96_271;
wire [0:0] comp_A994_365;
wire [0:0] comp_A999991_372;
wire [0:0] comp_A99999_168;
wire [0:0] comp_A95_430;
wire [0:0] comp_A8_398;
wire [0:0] comp_A994_484;
wire [0:0] comp_A999997_1009;
wire [0:0] comp_A3_415;
wire [0:0] comp_A97_174;
wire [0:0] comp_A997_549;
wire [0:0] comp_A999996_427;
wire [0:0] comp_A3_381;
wire [0:0] comp_A997_496;
wire [0:0] comp_A995_61;
wire [0:0] comp_A99_15;
wire [0:0] comp_A99_18;
wire [0:0] comp_A992_721;
wire [0:0] comp_A6_474;
wire [0:0] comp_A95_345;
wire [0:0] comp_A2_860;
wire [0:0] comp_A9_853;
wire [0:0] comp_A93_136;
wire [0:0] comp_A991_746;
wire [0:0] comp_A2_320;
wire [0:0] comp_A97_182;
wire [0:0] comp_A91_383;
wire [0:0] comp_A6_485;
wire [0:0] comp_A99995_471;
wire [0:0] comp_A93_516;
wire [0:0] comp_A99992_501;
wire [0:0] comp_A2_920;
wire [0:0] comp_A9991_961;
wire [0:0] comp_A999996_360;
wire [0:0] comp_A996_350;
wire [0:0] comp_A991_868;
wire [0:0] comp_A992_266;
wire [0:0] comp_A95_312;
wire [0:0] comp_A96_171;
wire [0:0] comp_A98_61;
wire [0:0] comp_A9994_693;
wire [0:0] comp_A994_378;
wire [0:0] comp_A99991_182;
wire [0:0] comp_A8_718;
wire [0:0] comp_A3_428;
wire [0:0] comp_A99996_862;
wire [0:0] comp_A9993_327;
wire [0:0] comp_A995_537;
wire [0:0] comp_A9_832;
wire [0:0] comp_A6_442;
wire [0:0] comp_A999996_428;
wire [0:0] comp_A94_58;
wire [0:0] comp_A997_521;
wire [0:0] comp_A996_360;
wire [0:0] comp_A99992_503;
wire [0:0] comp_A999994_457;
wire [0:0] comp_A99992_710;
wire [0:0] comp_A99991_366;
wire [0:0] comp_A993_286;
wire [0:0] comp_A999_567;
wire [0:0] comp_A99996_858;
wire [0:0] comp_A5_316;
wire [0:0] comp_A995_299;
wire [0:0] comp_A991_852;
wire [0:0] comp_A94_49;
wire [0:0] comp_A9992_105;
wire [0:0] comp_A92_247;
wire [0:0] comp_A98_68;
wire [0:0] comp_A99995_519;
wire [0:0] comp_A92_989;
wire [0:0] comp_A3_285;
wire [0:0] comp_A94_42;
wire [0:0] comp_A97_400;
wire [0:0] comp_A3_209;
wire [0:0] comp_A8_381;
wire [0:0] comp_A99_19;
wire [0:0] comp_A999997_1011;
wire [0:0] comp_A92_815;
wire [0:0] comp_A94_33;
wire [0:0] comp_A9991_937;
wire [0:0] comp_A998_499;
wire [0:0] comp_A1_554;
wire [0:0] comp_A999994_662;
wire [0:0] comp_A5_562;
wire [0:0] comp_A9997_669;
wire [0:0] comp_A997_477;
wire [0:0] comp_A9991_973;
wire [0:0] comp_A9999_248;
wire [0:0] comp_A996_245;
wire [0:0] comp_A98_1019;
wire [0:0] comp_A3_112;
wire [0:0] comp_A994_355;
wire [0:0] comp_A993_548;
wire [0:0] comp_A9991_817;
wire [0:0] comp_A92_246;
wire [0:0] comp_A3_27;
wire [0:0] comp_A8_810;
wire [0:0] comp_A99994_682;
wire [0:0] comp_A993_612;
wire [0:0] comp_A9992_99;
wire [0:0] comp_A9996_610;
wire [0:0] comp_A997_620;
wire [0:0] comp_A994_477;
wire [0:0] comp_A9999_293;
wire [0:0] comp_A8_404;
wire [0:0] comp_A996_318;
wire [0:0] comp_A95_274;
wire [0:0] comp_A1_601;
wire [0:0] comp_A92_562;
wire [0:0] comp_A99997_252;
wire [0:0] comp_A9996_694;
wire [0:0] comp_A3_305;
wire [0:0] comp_A997_334;
wire [0:0] comp_A999994_507;
wire [0:0] comp_A99993_647;
wire [0:0] comp_A992_308;
wire [0:0] comp_A99992_810;
wire [0:0] comp_A9993_652;
wire [0:0] comp_A997_403;
wire [0:0] comp_A93_651;
wire [0:0] comp_A999991_306;
wire [0:0] comp_A991_720;
wire [0:0] comp_A9992_107;
wire [0:0] comp_A9_851;
wire [0:0] comp_A9992_103;
wire [0:0] comp_A2_869;
wire [0:0] comp_A997_578;
wire [0:0] comp_A998_302;
wire [0:0] comp_A99991_660;
wire [0:0] comp_A6_644;
wire [0:0] comp_A2_285;
wire [0:0] comp_A995_202;
wire [0:0] comp_A8_818;
wire [0:0] comp_A999995_1012;
wire [0:0] comp_A997_956;
wire [0:0] comp_A999992_388;
wire [0:0] comp_A93_687;
wire [0:0] comp_A999995_1008;
wire [0:0] comp_A996_292;
wire [0:0] comp_A991_250;
wire [0:0] comp_A95_354;
wire [0:0] comp_A9994_711;
wire [0:0] comp_A9994_295;
wire [0:0] comp_A5_505;
wire [0:0] comp_A94_35;
wire [0:0] comp_A999994_547;
wire [0:0] comp_A9993_685;
wire [0:0] comp_A93_718;
wire [0:0] comp_A9991_956;
wire [0:0] comp_A993_484;
wire [0:0] comp_A1_708;
wire [0:0] comp_A9991_990;
wire [0:0] comp_A3_283;
wire [0:0] comp_A998_641;
wire [0:0] comp_A92_377;
wire [0:0] comp_A99994_383;
wire [0:0] comp_A999992_484;
wire [0:0] comp_A9_160;
wire [0:0] comp_A997_422;
wire [0:0] comp_A2_862;
wire [0:0] comp_A96_180;
wire [0:0] comp_A99997_843;
wire [0:0] comp_A9994_704;
wire [0:0] comp_A98_240;
wire [0:0] comp_A3_992;
wire [0:0] comp_A9994_881;
wire [0:0] comp_A2_827;
wire [0:0] comp_A999997_1012;
wire [0:0] comp_A994_549;
wire [0:0] comp_A97_171;
wire [0:0] comp_A9993_313;
wire [0:0] comp_A4_545;
wire [0:0] comp_A996_200;
wire [0:0] comp_A3_247;
wire [0:0] comp_A995_185;
wire [0:0] comp_A998_559;
wire [0:0] comp_A9999_767;
wire [0:0] comp_A99996_551;
wire [0:0] comp_A6_701;
wire [0:0] comp_A992_817;
wire [0:0] comp_A93_115;
wire [0:0] comp_A9991_962;
wire [0:0] comp_A99993_596;
wire [0:0] comp_A93_98;
wire [0:0] comp_A99994_807;
wire [0:0] comp_A96_264;
wire [0:0] comp_A92_500;
wire [0:0] comp_A9996_693;
wire [0:0] comp_A99993_630;
wire [0:0] comp_A99996_513;
wire [0:0] comp_A997_451;
wire [0:0] comp_A9992_161;
wire [0:0] comp_A2_114;
wire [0:0] comp_A995_493;
wire [0:0] comp_A99996_188;
wire [0:0] comp_A3_116;
wire [0:0] comp_A99996_839;
wire [0:0] comp_A2_9;
wire [0:0] comp_A93_544;
wire [0:0] comp_A3_812;
wire [0:0] comp_A997_373;
wire [0:0] comp_A99999_423;
wire [0:0] comp_A9991_955;
wire [0:0] comp_A9998_906;
wire [0:0] comp_A999996_461;
wire [0:0] comp_A999_585;
wire [0:0] comp_A5_753;
wire [0:0] comp_A99993_51;
wire [0:0] comp_A92_255;
wire [0:0] comp_A7_856;
wire [0:0] comp_A9_829;
wire [0:0] comp_A99995_559;
wire [0:0] comp_A2_33;
wire [0:0] comp_A99999_545;
wire [0:0] comp_A9992_436;
wire [0:0] comp_A997_666;
wire [0:0] comp_A94_37;
wire [0:0] comp_A9991_1011;
wire [0:0] comp_A99991_408;
wire [0:0] comp_A996_343;
wire [0:0] comp_A9999_560;
wire [0:0] comp_A996_263;
wire [0:0] comp_A9996_763;
wire [0:0] comp_A99992_660;
wire [0:0] comp_A1_642;
wire [0:0] comp_A9999_419;
wire [0:0] comp_A7_643;
wire [0:0] comp_A99992_736;
wire [0:0] comp_A9_61;
wire [0:0] comp_A6_394;
wire [0:0] comp_A99999_406;
wire [0:0] comp_A3_565;
wire [0:0] comp_A997_381;
wire [0:0] comp_A99992_538;
wire [0:0] comp_A99994_755;
wire [0:0] comp_A8_484;
wire [0:0] comp_A99992_655;
wire [0:0] comp_A991_451;
wire [0:0] comp_A99995_531;
wire [0:0] comp_A3_386;
wire [0:0] comp_A9998_389;
wire [0:0] comp_A994_390;
wire [0:0] comp_A97_201;
wire [0:0] comp_A3_750;
wire [0:0] comp_A995_34;
wire [0:0] comp_A994_677;
wire [0:0] comp_A93_720;
wire [0:0] comp_A99997_149;
wire [0:0] comp_A3_588;
wire [0:0] comp_A98_120;
wire [0:0] comp_A9_151;
wire [0:0] comp_A996_244;
wire [0:0] comp_A9999_786;
wire [0:0] comp_A99992_744;
wire [0:0] comp_A97_968;
wire [0:0] comp_A9993_626;
wire [0:0] comp_A99998_187;
wire [0:0] comp_A99994_612;
wire [0:0] comp_A9991_982;
wire [0:0] comp_A2_918;
wire [0:0] comp_A996_304;
wire [0:0] comp_A99_5;
wire [0:0] comp_A9991_693;
wire [0:0] comp_A99_21;
wire [0:0] comp_A9991_931;
wire [0:0] comp_A3_103;
wire [0:0] comp_A998_676;
wire [0:0] comp_A9_486;
wire [0:0] comp_A92_528;
wire [0:0] comp_A7_460;
wire [0:0] comp_A999994_411;
wire [0:0] comp_A93_722;
wire [0:0] comp_A98_153;
wire [0:0] comp_A996_231;
wire [0:0] comp_A999_516;
wire [0:0] comp_A991_373;
wire [0:0] comp_A9993_658;
wire [0:0] comp_A999992_474;
wire [0:0] comp_A999995_1014;
wire [0:0] comp_A9995_441;
wire [0:0] comp_A996_327;
wire [0:0] comp_A1_684;
wire [0:0] comp_A99999_443;
wire [0:0] comp_A9996_623;
wire [0:0] comp_A9_150;
wire [0:0] comp_A997_713;
wire [0:0] comp_A9991_965;
wire [0:0] comp_A999992_432;
wire [0:0] comp_A999996_726;
wire [0:0] comp_A993_258;
wire [0:0] comp_A8_335;
wire [0:0] comp_A999_656;
wire [0:0] comp_A991_735;
wire [0:0] comp_A996_203;
wire [0:0] comp_A93_546;
wire [0:0] comp_A99996_508;
wire [0:0] comp_A99996_263;
wire [0:0] comp_A9996_431;
wire [0:0] comp_A96_22;
wire [0:0] comp_A94_30;
wire [0:0] comp_A999_711;
wire [0:0] comp_A9_840;
wire [0:0] comp_A91_210;
wire [0:0] comp_A9997_587;
wire [0:0] comp_A2_713;
wire [0:0] comp_A999996_685;
wire [0:0] comp_A2_844;
wire [0:0] comp_A997_399;
wire [0:0] comp_A9993_561;
wire [0:0] comp_A991_391;
wire [0:0] comp_A6_286;
wire [0:0] comp_A99992_711;
wire [0:0] comp_A9991_921;
wire [0:0] comp_A3_55;
wire [0:0] comp_A9_157;
wire [0:0] comp_A8_657;
wire [0:0] comp_A99994_586;
wire [0:0] comp_A991_797;
wire [0:0] comp_A997_394;
wire [0:0] comp_A96_766;
wire [0:0] comp_A9993_581;
wire [0:0] comp_A9998_661;
wire [0:0] comp_A99993_699;
wire [0:0] comp_A9996_707;
wire [0:0] comp_A99997_955;
wire [0:0] comp_A991_647;
wire [0:0] comp_A996_185;
wire [0:0] comp_A999992_536;
wire [0:0] comp_A93_92;
wire [0:0] comp_A1_581;
wire [0:0] comp_A991_486;
wire [0:0] comp_A993_621;
wire [0:0] comp_A999992_339;
wire [0:0] comp_A7_767;
wire [0:0] comp_A99993_85;
wire [0:0] comp_A92_574;
wire [0:0] comp_A3_867;
wire [0:0] comp_A98_270;
wire [0:0] comp_A93_119;
wire [0:0] comp_A992_234;
wire [0:0] comp_A92_992;
wire [0:0] comp_A991_644;
wire [0:0] comp_A3_662;
wire [0:0] comp_A996_311;
wire [0:0] comp_A994_457;
wire [0:0] comp_A9993_539;
wire [0:0] comp_A99997_946;
wire [0:0] comp_A997_299;
wire [0:0] comp_A99992_670;
wire [0:0] comp_A94_32;
wire [0:0] comp_A1_741;
wire [0:0] comp_A994_524;
wire [0:0] comp_A9997_340;
wire [0:0] comp_A997_696;
wire [0:0] comp_A99994_727;
wire [0:0] comp_A994_644;
wire [0:0] comp_A996_369;
wire [0:0] comp_A9991_995;
wire [0:0] comp_A5_492;
wire [0:0] comp_A998_230;
wire [0:0] comp_A93_532;
wire [0:0] comp_A999_337;
wire [0:0] comp_A95_388;
wire [0:0] comp_A3_127;
wire [0:0] comp_A6_452;
wire [0:0] comp_A4_332;
wire [0:0] comp_A999996_581;
wire [0:0] comp_A8_875;
wire [0:0] comp_A97_207;
wire [0:0] comp_A9993_671;
wire [0:0] comp_A9999_59;
wire [0:0] comp_A991_777;
wire [0:0] comp_A9991_699;
COMPS INST_COMP(
reg_A1, reg_A2, reg_A3, reg_A4, reg_A5, reg_A6, reg_A7, reg_A8, reg_A9, reg_A91, reg_A92, reg_A93, reg_A94, reg_A95, reg_A96, reg_A97, reg_A98, reg_A99, reg_A991, reg_A992, reg_A993, reg_A994, reg_A995, reg_A996, reg_A997, reg_A998, reg_A999, reg_A9991, reg_A9992, reg_A9993, reg_A9994, reg_A9995, reg_A9996, reg_A9997, reg_A9998, reg_A9999, reg_A99991, reg_A99992, reg_A99993, reg_A99994, reg_A99995, reg_A99996, reg_A99997, reg_A99998, reg_A99999, reg_A999991, reg_A999992, reg_A999993, reg_A999994, reg_A999995, reg_A999996, reg_A999997, comp_A1_649, comp_A2_29, comp_A3_322, comp_A4_504, comp_A5_495, comp_A6_624, comp_A7_593, comp_A1_220, comp_A4_472, comp_A8_701, comp_A9_178, comp_A91_362, comp_A92_263, comp_A93_529, comp_A94_40, comp_A7_795, comp_A95_118, comp_A3_541, comp_A8_90, comp_A96_11, comp_A97_193, comp_A98_202, comp_A99_14, comp_A2_830, comp_A991_288, comp_A992_452, comp_A95_373, comp_A8_777, comp_A93_537, comp_A99_11, comp_A95_383, comp_A993_454, comp_A992_774, comp_A994_302, comp_A995_87, comp_A98_143, comp_A996_348, comp_A997_750, comp_A1_884, comp_A997_360, comp_A998_765, comp_A8_726, comp_A999_643, comp_A3_526, comp_A7_455, comp_A9991_920, comp_A3_300, comp_A92_262, comp_A9992_183, comp_A991_737, comp_A97_140, comp_A9991_923, comp_A96_873, comp_A9993_513, comp_A4_515, comp_A9994_577, comp_A94_46, comp_A7_341, comp_A3_687, comp_A9995_483, comp_A9996_660, comp_A9997_526, comp_A9991_943, comp_A7_561, comp_A993_276, comp_A9998_478, comp_A92_975, comp_A1_727, comp_A7_583, comp_A995_79, comp_A97_173, comp_A993_665, comp_A9999_801, comp_A3_536, comp_A999_620, comp_A994_700, comp_A99991_242, comp_A994_712, comp_A99992_806, comp_A9997_570, comp_A99993_119, comp_A6_670, comp_A994_338, comp_A6_635, comp_A9994_627, comp_A1_881, comp_A4_490, comp_A92_264, comp_A2_839, comp_A991_760, comp_A993_680, comp_A99994_810, comp_A98_974, comp_A4_350, comp_A1_738, comp_A997_319, comp_A7_411, comp_A4_400, comp_A9992_93, comp_A99994_781, comp_A93_726, comp_A9998_769, comp_A7_415, comp_A9991_972, comp_A993_608, comp_A3_284, comp_A9995_876, comp_A9_859, comp_A9992_129, comp_A3_102, comp_A3_79, comp_A9993_585, comp_A3_124, comp_A91_239, comp_A93_116, comp_A9_811, comp_A3_757, comp_A99991_336, comp_A98_66, comp_A99995_631, comp_A999_732, comp_A9996_244, comp_A995_167, comp_A98_171, comp_A3_981, comp_A9_827, comp_A9992_357, comp_A4_739, comp_A2_876, comp_A99996_412, comp_A9996_202, comp_A9993_525, comp_A7_666, comp_A92_519, comp_A99994_745, comp_A998_448, comp_A9997_490, comp_A9996_448, comp_A997_332, comp_A4_495, comp_A94_29, comp_A7_919, comp_A99997_247, comp_A993_764, comp_A9991_914, comp_A96_609, comp_A9999_832, comp_A99998_189, comp_A996_296, comp_A99999_409, comp_A99994_713, comp_A993_839, comp_A99997_833, comp_A5_327, comp_A2_894, comp_A3_587, comp_A93_629, comp_A999991_302, comp_A99997_824, comp_A9_155, comp_A5_170, comp_A97_991, comp_A995_114, comp_A5_586, comp_A98_162, comp_A991_728, comp_A9996_782, comp_A99992_505, comp_A9995_733, comp_A9991_1016, comp_A9_152, comp_A5_126, comp_A999992_426, comp_A9_784, comp_A999992_487, comp_A92_504, comp_A9994_769, comp_A95_435, comp_A999992_569, comp_A1_652, comp_A991_268, comp_A99997_799, comp_A992_599, comp_A99991_539, comp_A98_147, comp_A7_591, comp_A997_589, comp_A97_124, comp_A996_225, comp_A97_121, comp_A99995_671, comp_A9998_723, comp_A999993_9, comp_A996_92, comp_A996_222, comp_A9999_756, comp_A95_203, comp_A997_838, comp_A5_478, comp_A99997_254, comp_A99991_618, comp_A91_963, comp_A9994_288, comp_A9991_935, comp_A99997_931, comp_A98_151, comp_A4_486, comp_A3_232, comp_A9995_839, comp_A7_592, comp_A3_286, comp_A99999_486, comp_A9991_932, comp_A996_372, comp_A9_156, comp_A7_804, comp_A6_255, comp_A99991_344, comp_A8_757, comp_A993_555, comp_A999994_442, comp_A99992_671, comp_A991_479, comp_A97_610, comp_A999991_570, comp_A9_816, comp_A3_80, comp_A8_822, comp_A998_424, comp_A999993_8, comp_A9992_421, comp_A99999_549, comp_A9993_307, comp_A9996_562, comp_A996_271, comp_A992_400, comp_A94_31, comp_A99_8, comp_A3_54, comp_A2_872, comp_A92_972, comp_A3_272, comp_A999995_1015, comp_A7_605, comp_A9993_295, comp_A991_531, comp_A993_317, comp_A991_869, comp_A94_50, comp_A99994_178, comp_A8_786, comp_A3_407, comp_A6_722, comp_A99999_735, comp_A92_259, comp_A999996_390, comp_A2_901, comp_A992_675, comp_A9_821, comp_A92_503, comp_A8_536, comp_A2_124, comp_A92_250, comp_A95_497, comp_A6_406, comp_A9991_948, comp_A9999_819, comp_A3_535, comp_A998_805, comp_A92_995, comp_A9996_600, comp_A6_606, comp_A996_353, comp_A99994_600, comp_A99991_286, comp_A996_340, comp_A998_414, comp_A996_331, comp_A994_640, comp_A999_714, comp_A3_233, comp_A9_805, comp_A8_540, comp_A99996_575, comp_A993_982, comp_A9993_530, comp_A994_475, comp_A996_332, comp_A4_484, comp_A98_325, comp_A993_659, comp_A2_602, comp_A92_505, comp_A99999_58, comp_A9992_123, comp_A999992_527, comp_A9996_758, comp_A997_428, comp_A3_515, comp_A992_389, comp_A93_513, comp_A99999_558, comp_A9992_429, comp_A993_440, comp_A99996_766, comp_A999991_485, comp_A9991_1009, comp_A99999_594, comp_A993_492, comp_A96_754, comp_A993_321, comp_A999_712, comp_A997_421, comp_A9999_805, comp_A995_343, comp_A9996_570, comp_A5_653, comp_A4_445, comp_A99995_511, comp_A99991_185, comp_A99999_517, comp_A8_334, comp_A9996_737, comp_A9_845, comp_A997_339, comp_A997_243, comp_A993_683, comp_A994_543, comp_A99_13, comp_A2_22, comp_A96_818, comp_A3_350, comp_A992_528, comp_A96_271, comp_A994_365, comp_A999991_372, comp_A99999_168, comp_A95_430, comp_A8_398, comp_A994_484, comp_A999997_1009, comp_A3_415, comp_A97_174, comp_A997_549, comp_A999996_427, comp_A3_381, comp_A997_496, comp_A995_61, comp_A99_15, comp_A99_18, comp_A992_721, comp_A6_474, comp_A95_345, comp_A2_860, comp_A9_853, comp_A93_136, comp_A991_746, comp_A2_320, comp_A97_182, comp_A91_383, comp_A6_485, comp_A99995_471, comp_A93_516, comp_A99992_501, comp_A2_920, comp_A9991_961, comp_A999996_360, comp_A996_350, comp_A991_868, comp_A992_266, comp_A95_312, comp_A96_171, comp_A98_61, comp_A9994_693, comp_A994_378, comp_A99991_182, comp_A8_718, comp_A3_428, comp_A99996_862, comp_A9993_327, comp_A995_537, comp_A9_832, comp_A6_442, comp_A999996_428, comp_A94_58, comp_A997_521, comp_A996_360, comp_A99992_503, comp_A999994_457, comp_A99992_710, comp_A99991_366, comp_A993_286, comp_A999_567, comp_A99996_858, comp_A5_316, comp_A995_299, comp_A991_852, comp_A94_49, comp_A9992_105, comp_A92_247, comp_A98_68, comp_A99995_519, comp_A92_989, comp_A3_285, comp_A94_42, comp_A97_400, comp_A3_209, comp_A8_381, comp_A99_19, comp_A999997_1011, comp_A92_815, comp_A94_33, comp_A9991_937, comp_A998_499, comp_A1_554, comp_A999994_662, comp_A5_562, comp_A9997_669, comp_A997_477, comp_A9991_973, comp_A9999_248, comp_A996_245, comp_A98_1019, comp_A3_112, comp_A994_355, comp_A993_548, comp_A9991_817, comp_A92_246, comp_A3_27, comp_A8_810, comp_A99994_682, comp_A993_612, comp_A9992_99, comp_A9996_610, comp_A997_620, comp_A994_477, comp_A9999_293, comp_A8_404, comp_A996_318, comp_A95_274, comp_A1_601, comp_A92_562, comp_A99997_252, comp_A9996_694, comp_A3_305, comp_A997_334, comp_A999994_507, comp_A99993_647, comp_A992_308, comp_A99992_810, comp_A9993_652, comp_A997_403, comp_A93_651, comp_A999991_306, comp_A991_720, comp_A9992_107, comp_A9_851, comp_A9992_103, comp_A2_869, comp_A997_578, comp_A998_302, comp_A99991_660, comp_A6_644, comp_A2_285, comp_A995_202, comp_A8_818, comp_A999995_1012, comp_A997_956, comp_A999992_388, comp_A93_687, comp_A999995_1008, comp_A996_292, comp_A991_250, comp_A95_354, comp_A9994_711, comp_A9994_295, comp_A5_505, comp_A94_35, comp_A999994_547, comp_A9993_685, comp_A93_718, comp_A9991_956, comp_A993_484, comp_A1_708, comp_A9991_990, comp_A3_283, comp_A998_641, comp_A92_377, comp_A99994_383, comp_A999992_484, comp_A9_160, comp_A997_422, comp_A2_862, comp_A96_180, comp_A99997_843, comp_A9994_704, comp_A98_240, comp_A3_992, comp_A9994_881, comp_A2_827, comp_A999997_1012, comp_A994_549, comp_A97_171, comp_A9993_313, comp_A4_545, comp_A996_200, comp_A3_247, comp_A995_185, comp_A998_559, comp_A9999_767, comp_A99996_551, comp_A6_701, comp_A992_817, comp_A93_115, comp_A9991_962, comp_A99993_596, comp_A93_98, comp_A99994_807, comp_A96_264, comp_A92_500, comp_A9996_693, comp_A99993_630, comp_A99996_513, comp_A997_451, comp_A9992_161, comp_A2_114, comp_A995_493, comp_A99996_188, comp_A3_116, comp_A99996_839, comp_A2_9, comp_A93_544, comp_A3_812, comp_A997_373, comp_A99999_423, comp_A9991_955, comp_A9998_906, comp_A999996_461, comp_A999_585, comp_A5_753, comp_A99993_51, comp_A92_255, comp_A7_856, comp_A9_829, comp_A99995_559, comp_A2_33, comp_A99999_545, comp_A9992_436, comp_A997_666, comp_A94_37, comp_A9991_1011, comp_A99991_408, comp_A996_343, comp_A9999_560, comp_A996_263, comp_A9996_763, comp_A99992_660, comp_A1_642, comp_A9999_419, comp_A7_643, comp_A99992_736, comp_A9_61, comp_A6_394, comp_A99999_406, comp_A3_565, comp_A997_381, comp_A99992_538, comp_A99994_755, comp_A8_484, comp_A99992_655, comp_A991_451, comp_A99995_531, comp_A3_386, comp_A9998_389, comp_A994_390, comp_A97_201, comp_A3_750, comp_A995_34, comp_A994_677, comp_A93_720, comp_A99997_149, comp_A3_588, comp_A98_120, comp_A9_151, comp_A996_244, comp_A9999_786, comp_A99992_744, comp_A97_968, comp_A9993_626, comp_A99998_187, comp_A99994_612, comp_A9991_982, comp_A2_918, comp_A996_304, comp_A99_5, comp_A9991_693, comp_A99_21, comp_A9991_931, comp_A3_103, comp_A998_676, comp_A9_486, comp_A92_528, comp_A7_460, comp_A999994_411, comp_A93_722, comp_A98_153, comp_A996_231, comp_A999_516, comp_A991_373, comp_A9993_658, comp_A999992_474, comp_A999995_1014, comp_A9995_441, comp_A996_327, comp_A1_684, comp_A99999_443, comp_A9996_623, comp_A9_150, comp_A997_713, comp_A9991_965, comp_A999992_432, comp_A999996_726, comp_A993_258, comp_A8_335, comp_A999_656, comp_A991_735, comp_A996_203, comp_A93_546, comp_A99996_508, comp_A99996_263, comp_A9996_431, comp_A96_22, comp_A94_30, comp_A999_711, comp_A9_840, comp_A91_210, comp_A9997_587, comp_A2_713, comp_A999996_685, comp_A2_844, comp_A997_399, comp_A9993_561, comp_A991_391, comp_A6_286, comp_A99992_711, comp_A9991_921, comp_A3_55, comp_A9_157, comp_A8_657, comp_A99994_586, comp_A991_797, comp_A997_394, comp_A96_766, comp_A9993_581, comp_A9998_661, comp_A99993_699, comp_A9996_707, comp_A99997_955, comp_A991_647, comp_A996_185, comp_A999992_536, comp_A93_92, comp_A1_581, comp_A991_486, comp_A993_621, comp_A999992_339, comp_A7_767, comp_A99993_85, comp_A92_574, comp_A3_867, comp_A98_270, comp_A93_119, comp_A992_234, comp_A92_992, comp_A991_644, comp_A3_662, comp_A996_311, comp_A994_457, comp_A9993_539, comp_A99997_946, comp_A997_299, comp_A99992_670, comp_A94_32, comp_A1_741, comp_A994_524, comp_A9997_340, comp_A997_696, comp_A99994_727, comp_A994_644, comp_A996_369, comp_A9991_995, comp_A5_492, comp_A998_230, comp_A93_532, comp_A999_337, comp_A95_388, comp_A3_127, comp_A6_452, comp_A4_332, comp_A999996_581, comp_A8_875, comp_A97_207, comp_A9993_671, comp_A9999_59, comp_A991_777, comp_A9991_699
);

ANDS INST_ANDS(
comp_A1_649, comp_A2_29, comp_A3_322, comp_A4_504, comp_A5_495, comp_A6_624, comp_A7_593, comp_A1_220, comp_A4_472, comp_A8_701, comp_A9_178, comp_A91_362, comp_A92_263, comp_A93_529, comp_A94_40, comp_A7_795, comp_A95_118, comp_A3_541, comp_A8_90, comp_A96_11, comp_A97_193, comp_A98_202, comp_A99_14, comp_A2_830, comp_A991_288, comp_A992_452, comp_A95_373, comp_A8_777, comp_A93_537, comp_A99_11, comp_A95_383, comp_A993_454, comp_A992_774, comp_A994_302, comp_A995_87, comp_A98_143, comp_A996_348, comp_A997_750, comp_A1_884, comp_A997_360, comp_A998_765, comp_A8_726, comp_A999_643, comp_A3_526, comp_A7_455, comp_A9991_920, comp_A3_300, comp_A92_262, comp_A9992_183, comp_A991_737, comp_A97_140, comp_A9991_923, comp_A96_873, comp_A9993_513, comp_A4_515, comp_A9994_577, comp_A94_46, comp_A7_341, comp_A3_687, comp_A9995_483, comp_A9996_660, comp_A9997_526, comp_A9991_943, comp_A7_561, comp_A993_276, comp_A9998_478, comp_A92_975, comp_A1_727, comp_A7_583, comp_A995_79, comp_A97_173, comp_A993_665, comp_A9999_801, comp_A3_536, comp_A999_620, comp_A994_700, comp_A99991_242, comp_A994_712, comp_A99992_806, comp_A9997_570, comp_A99993_119, comp_A6_670, comp_A994_338, comp_A6_635, comp_A9994_627, comp_A1_881, comp_A4_490, comp_A92_264, comp_A2_839, comp_A991_760, comp_A993_680, comp_A99994_810, comp_A98_974, comp_A4_350, comp_A1_738, comp_A997_319, comp_A7_411, comp_A4_400, comp_A9992_93, comp_A99994_781, comp_A93_726, comp_A9998_769, comp_A7_415, comp_A9991_972, comp_A993_608, comp_A3_284, comp_A9995_876, comp_A9_859, comp_A9992_129, comp_A3_102, comp_A3_79, comp_A9993_585, comp_A3_124, comp_A91_239, comp_A93_116, comp_A9_811, comp_A3_757, comp_A99991_336, comp_A98_66, comp_A99995_631, comp_A999_732, comp_A9996_244, comp_A995_167, comp_A98_171, comp_A3_981, comp_A9_827, comp_A9992_357, comp_A4_739, comp_A2_876, comp_A99996_412, comp_A9996_202, comp_A9993_525, comp_A7_666, comp_A92_519, comp_A99994_745, comp_A998_448, comp_A9997_490, comp_A9996_448, comp_A997_332, comp_A4_495, comp_A94_29, comp_A7_919, comp_A99997_247, comp_A993_764, comp_A9991_914, comp_A96_609, comp_A9999_832, comp_A99998_189, comp_A996_296, comp_A99999_409, comp_A99994_713, comp_A993_839, comp_A99997_833, comp_A5_327, comp_A2_894, comp_A3_587, comp_A93_629, comp_A999991_302, comp_A99997_824, comp_A9_155, comp_A5_170, comp_A97_991, comp_A995_114, comp_A5_586, comp_A98_162, comp_A991_728, comp_A9996_782, comp_A99992_505, comp_A9995_733, comp_A9991_1016, comp_A9_152, comp_A5_126, comp_A999992_426, comp_A9_784, comp_A999992_487, comp_A92_504, comp_A9994_769, comp_A95_435, comp_A999992_569, comp_A1_652, comp_A991_268, comp_A99997_799, comp_A992_599, comp_A99991_539, comp_A98_147, comp_A7_591, comp_A997_589, comp_A97_124, comp_A996_225, comp_A97_121, comp_A99995_671, comp_A9998_723, comp_A999993_9, comp_A996_92, comp_A996_222, comp_A9999_756, comp_A95_203, comp_A997_838, comp_A5_478, comp_A99997_254, comp_A99991_618, comp_A91_963, comp_A9994_288, comp_A9991_935, comp_A99997_931, comp_A98_151, comp_A4_486, comp_A3_232, comp_A9995_839, comp_A7_592, comp_A3_286, comp_A99999_486, comp_A9991_932, comp_A996_372, comp_A9_156, comp_A7_804, comp_A6_255, comp_A99991_344, comp_A8_757, comp_A993_555, comp_A999994_442, comp_A99992_671, comp_A991_479, comp_A97_610, comp_A999991_570, comp_A9_816, comp_A3_80, comp_A8_822, comp_A998_424, comp_A999993_8, comp_A9992_421, comp_A99999_549, comp_A9993_307, comp_A9996_562, comp_A996_271, comp_A992_400, comp_A94_31, comp_A99_8, comp_A3_54, comp_A2_872, comp_A92_972, comp_A3_272, comp_A999995_1015, comp_A7_605, comp_A9993_295, comp_A991_531, comp_A993_317, comp_A991_869, comp_A94_50, comp_A99994_178, comp_A8_786, comp_A3_407, comp_A6_722, comp_A99999_735, comp_A92_259, comp_A999996_390, comp_A2_901, comp_A992_675, comp_A9_821, comp_A92_503, comp_A8_536, comp_A2_124, comp_A92_250, comp_A95_497, comp_A6_406, comp_A9991_948, comp_A9999_819, comp_A3_535, comp_A998_805, comp_A92_995, comp_A9996_600, comp_A6_606, comp_A996_353, comp_A99994_600, comp_A99991_286, comp_A996_340, comp_A998_414, comp_A996_331, comp_A994_640, comp_A999_714, comp_A3_233, comp_A9_805, comp_A8_540, comp_A99996_575, comp_A993_982, comp_A9993_530, comp_A994_475, comp_A996_332, comp_A4_484, comp_A98_325, comp_A993_659, comp_A2_602, comp_A92_505, comp_A99999_58, comp_A9992_123, comp_A999992_527, comp_A9996_758, comp_A997_428, comp_A3_515, comp_A992_389, comp_A93_513, comp_A99999_558, comp_A9992_429, comp_A993_440, comp_A99996_766, comp_A999991_485, comp_A9991_1009, comp_A99999_594, comp_A993_492, comp_A96_754, comp_A993_321, comp_A999_712, comp_A997_421, comp_A9999_805, comp_A995_343, comp_A9996_570, comp_A5_653, comp_A4_445, comp_A99995_511, comp_A99991_185, comp_A99999_517, comp_A8_334, comp_A9996_737, comp_A9_845, comp_A997_339, comp_A997_243, comp_A993_683, comp_A994_543, comp_A99_13, comp_A2_22, comp_A96_818, comp_A3_350, comp_A992_528, comp_A96_271, comp_A994_365, comp_A999991_372, comp_A99999_168, comp_A95_430, comp_A8_398, comp_A994_484, comp_A999997_1009, comp_A3_415, comp_A97_174, comp_A997_549, comp_A999996_427, comp_A3_381, comp_A997_496, comp_A995_61, comp_A99_15, comp_A99_18, comp_A992_721, comp_A6_474, comp_A95_345, comp_A2_860, comp_A9_853, comp_A93_136, comp_A991_746, comp_A2_320, comp_A97_182, comp_A91_383, comp_A6_485, comp_A99995_471, comp_A93_516, comp_A99992_501, comp_A2_920, comp_A9991_961, comp_A999996_360, comp_A996_350, comp_A991_868, comp_A992_266, comp_A95_312, comp_A96_171, comp_A98_61, comp_A9994_693, comp_A994_378, comp_A99991_182, comp_A8_718, comp_A3_428, comp_A99996_862, comp_A9993_327, comp_A995_537, comp_A9_832, comp_A6_442, comp_A999996_428, comp_A94_58, comp_A997_521, comp_A996_360, comp_A99992_503, comp_A999994_457, comp_A99992_710, comp_A99991_366, comp_A993_286, comp_A999_567, comp_A99996_858, comp_A5_316, comp_A995_299, comp_A991_852, comp_A94_49, comp_A9992_105, comp_A92_247, comp_A98_68, comp_A99995_519, comp_A92_989, comp_A3_285, comp_A94_42, comp_A97_400, comp_A3_209, comp_A8_381, comp_A99_19, comp_A999997_1011, comp_A92_815, comp_A94_33, comp_A9991_937, comp_A998_499, comp_A1_554, comp_A999994_662, comp_A5_562, comp_A9997_669, comp_A997_477, comp_A9991_973, comp_A9999_248, comp_A996_245, comp_A98_1019, comp_A3_112, comp_A994_355, comp_A993_548, comp_A9991_817, comp_A92_246, comp_A3_27, comp_A8_810, comp_A99994_682, comp_A993_612, comp_A9992_99, comp_A9996_610, comp_A997_620, comp_A994_477, comp_A9999_293, comp_A8_404, comp_A996_318, comp_A95_274, comp_A1_601, comp_A92_562, comp_A99997_252, comp_A9996_694, comp_A3_305, comp_A997_334, comp_A999994_507, comp_A99993_647, comp_A992_308, comp_A99992_810, comp_A9993_652, comp_A997_403, comp_A93_651, comp_A999991_306, comp_A991_720, comp_A9992_107, comp_A9_851, comp_A9992_103, comp_A2_869, comp_A997_578, comp_A998_302, comp_A99991_660, comp_A6_644, comp_A2_285, comp_A995_202, comp_A8_818, comp_A999995_1012, comp_A997_956, comp_A999992_388, comp_A93_687, comp_A999995_1008, comp_A996_292, comp_A991_250, comp_A95_354, comp_A9994_711, comp_A9994_295, comp_A5_505, comp_A94_35, comp_A999994_547, comp_A9993_685, comp_A93_718, comp_A9991_956, comp_A993_484, comp_A1_708, comp_A9991_990, comp_A3_283, comp_A998_641, comp_A92_377, comp_A99994_383, comp_A999992_484, comp_A9_160, comp_A997_422, comp_A2_862, comp_A96_180, comp_A99997_843, comp_A9994_704, comp_A98_240, comp_A3_992, comp_A9994_881, comp_A2_827, comp_A999997_1012, comp_A994_549, comp_A97_171, comp_A9993_313, comp_A4_545, comp_A996_200, comp_A3_247, comp_A995_185, comp_A998_559, comp_A9999_767, comp_A99996_551, comp_A6_701, comp_A992_817, comp_A93_115, comp_A9991_962, comp_A99993_596, comp_A93_98, comp_A99994_807, comp_A96_264, comp_A92_500, comp_A9996_693, comp_A99993_630, comp_A99996_513, comp_A997_451, comp_A9992_161, comp_A2_114, comp_A995_493, comp_A99996_188, comp_A3_116, comp_A99996_839, comp_A2_9, comp_A93_544, comp_A3_812, comp_A997_373, comp_A99999_423, comp_A9991_955, comp_A9998_906, comp_A999996_461, comp_A999_585, comp_A5_753, comp_A99993_51, comp_A92_255, comp_A7_856, comp_A9_829, comp_A99995_559, comp_A2_33, comp_A99999_545, comp_A9992_436, comp_A997_666, comp_A94_37, comp_A9991_1011, comp_A99991_408, comp_A996_343, comp_A9999_560, comp_A996_263, comp_A9996_763, comp_A99992_660, comp_A1_642, comp_A9999_419, comp_A7_643, comp_A99992_736, comp_A9_61, comp_A6_394, comp_A99999_406, comp_A3_565, comp_A997_381, comp_A99992_538, comp_A99994_755, comp_A8_484, comp_A99992_655, comp_A991_451, comp_A99995_531, comp_A3_386, comp_A9998_389, comp_A994_390, comp_A97_201, comp_A3_750, comp_A995_34, comp_A994_677, comp_A93_720, comp_A99997_149, comp_A3_588, comp_A98_120, comp_A9_151, comp_A996_244, comp_A9999_786, comp_A99992_744, comp_A97_968, comp_A9993_626, comp_A99998_187, comp_A99994_612, comp_A9991_982, comp_A2_918, comp_A996_304, comp_A99_5, comp_A9991_693, comp_A99_21, comp_A9991_931, comp_A3_103, comp_A998_676, comp_A9_486, comp_A92_528, comp_A7_460, comp_A999994_411, comp_A93_722, comp_A98_153, comp_A996_231, comp_A999_516, comp_A991_373, comp_A9993_658, comp_A999992_474, comp_A999995_1014, comp_A9995_441, comp_A996_327, comp_A1_684, comp_A99999_443, comp_A9996_623, comp_A9_150, comp_A997_713, comp_A9991_965, comp_A999992_432, comp_A999996_726, comp_A993_258, comp_A8_335, comp_A999_656, comp_A991_735, comp_A996_203, comp_A93_546, comp_A99996_508, comp_A99996_263, comp_A9996_431, comp_A96_22, comp_A94_30, comp_A999_711, comp_A9_840, comp_A91_210, comp_A9997_587, comp_A2_713, comp_A999996_685, comp_A2_844, comp_A997_399, comp_A9993_561, comp_A991_391, comp_A6_286, comp_A99992_711, comp_A9991_921, comp_A3_55, comp_A9_157, comp_A8_657, comp_A99994_586, comp_A991_797, comp_A997_394, comp_A96_766, comp_A9993_581, comp_A9998_661, comp_A99993_699, comp_A9996_707, comp_A99997_955, comp_A991_647, comp_A996_185, comp_A999992_536, comp_A93_92, comp_A1_581, comp_A991_486, comp_A993_621, comp_A999992_339, comp_A7_767, comp_A99993_85, comp_A92_574, comp_A3_867, comp_A98_270, comp_A93_119, comp_A992_234, comp_A92_992, comp_A991_644, comp_A3_662, comp_A996_311, comp_A994_457, comp_A9993_539, comp_A99997_946, comp_A997_299, comp_A99992_670, comp_A94_32, comp_A1_741, comp_A994_524, comp_A9997_340, comp_A997_696, comp_A99994_727, comp_A994_644, comp_A996_369, comp_A9991_995, comp_A5_492, comp_A998_230, comp_A93_532, comp_A999_337, comp_A95_388, comp_A3_127, comp_A6_452, comp_A4_332, comp_A999996_581, comp_A8_875, comp_A97_207, comp_A9993_671, comp_A9999_59, comp_A991_777, comp_A9991_699, or_0, or_1, or_2, or_3, or_4, or_5, or_6, or_7, or_8, or_9, or_10, or_11, or_12, or_13, or_14, or_15, or_16, or_17, or_18, or_19, or_20, or_21, or_22, or_23, or_24
);

MAJ INST_MAJ(
or_0, or_1, or_2, or_3, or_4, or_5, or_6, or_7, or_8, or_9, or_10, or_11, or_12, or_13, or_14, or_15, or_16, or_17, or_18, or_19, or_20, or_21, or_22, or_23, or_24, reg_decision
);


	assign reg_A1 = A1;

	assign reg_A2 = A2;

	assign reg_A3 = A3;

	assign reg_A4 = A4;

	assign reg_A5 = A5;

	assign reg_A6 = A6;

	assign reg_A7 = A7;

	assign reg_A8 = A8;

	assign reg_A9 = A9;

	assign reg_A91 = A91;

	assign reg_A92 = A92;

	assign reg_A93 = A93;

	assign reg_A94 = A94;

	assign reg_A95 = A95;

	assign reg_A96 = A96;

	assign reg_A97 = A97;

	assign reg_A98 = A98;

	assign reg_A99 = A99;

	assign reg_A991 = A991;

	assign reg_A992 = A992;

	assign reg_A993 = A993;

	assign reg_A994 = A994;

	assign reg_A995 = A995;

	assign reg_A996 = A996;

	assign reg_A997 = A997;

	assign reg_A998 = A998;

	assign reg_A999 = A999;

	assign reg_A9991 = A9991;

	assign reg_A9992 = A9992;

	assign reg_A9993 = A9993;

	assign reg_A9994 = A9994;

	assign reg_A9995 = A9995;

	assign reg_A9996 = A9996;

	assign reg_A9997 = A9997;

	assign reg_A9998 = A9998;

	assign reg_A9999 = A9999;

	assign reg_A99991 = A99991;

	assign reg_A99992 = A99992;

	assign reg_A99993 = A99993;

	assign reg_A99994 = A99994;

	assign reg_A99995 = A99995;

	assign reg_A99996 = A99996;

	assign reg_A99997 = A99997;

	assign reg_A99998 = A99998;

	assign reg_A99999 = A99999;

	assign reg_A999991 = A999991;

	assign reg_A999992 = A999992;

	assign reg_A999993 = A999993;

	assign reg_A999994 = A999994;

	assign reg_A999995 = A999995;

	assign reg_A999996 = A999996;

	assign reg_A999997 = A999997;

	assign decision = reg_decision;

endmodule


module COMPS(
reg_A1, reg_A2, reg_A3, reg_A4, reg_A5, reg_A6, reg_A7, reg_A8, reg_A9, reg_A91, reg_A92, reg_A93, reg_A94, reg_A95, reg_A96, reg_A97, reg_A98, reg_A99, reg_A991, reg_A992, reg_A993, reg_A994, reg_A995, reg_A996, reg_A997, reg_A998, reg_A999, reg_A9991, reg_A9992, reg_A9993, reg_A9994, reg_A9995, reg_A9996, reg_A9997, reg_A9998, reg_A9999, reg_A99991, reg_A99992, reg_A99993, reg_A99994, reg_A99995, reg_A99996, reg_A99997, reg_A99998, reg_A99999, reg_A999991, reg_A999992, reg_A999993, reg_A999994, reg_A999995, reg_A999996, reg_A999997, comp_A1_649, comp_A2_29, comp_A3_322, comp_A4_504, comp_A5_495, comp_A6_624, comp_A7_593, comp_A1_220, comp_A4_472, comp_A8_701, comp_A9_178, comp_A91_362, comp_A92_263, comp_A93_529, comp_A94_40, comp_A7_795, comp_A95_118, comp_A3_541, comp_A8_90, comp_A96_11, comp_A97_193, comp_A98_202, comp_A99_14, comp_A2_830, comp_A991_288, comp_A992_452, comp_A95_373, comp_A8_777, comp_A93_537, comp_A99_11, comp_A95_383, comp_A993_454, comp_A992_774, comp_A994_302, comp_A995_87, comp_A98_143, comp_A996_348, comp_A997_750, comp_A1_884, comp_A997_360, comp_A998_765, comp_A8_726, comp_A999_643, comp_A3_526, comp_A7_455, comp_A9991_920, comp_A3_300, comp_A92_262, comp_A9992_183, comp_A991_737, comp_A97_140, comp_A9991_923, comp_A96_873, comp_A9993_513, comp_A4_515, comp_A9994_577, comp_A94_46, comp_A7_341, comp_A3_687, comp_A9995_483, comp_A9996_660, comp_A9997_526, comp_A9991_943, comp_A7_561, comp_A993_276, comp_A9998_478, comp_A92_975, comp_A1_727, comp_A7_583, comp_A995_79, comp_A97_173, comp_A993_665, comp_A9999_801, comp_A3_536, comp_A999_620, comp_A994_700, comp_A99991_242, comp_A994_712, comp_A99992_806, comp_A9997_570, comp_A99993_119, comp_A6_670, comp_A994_338, comp_A6_635, comp_A9994_627, comp_A1_881, comp_A4_490, comp_A92_264, comp_A2_839, comp_A991_760, comp_A993_680, comp_A99994_810, comp_A98_974, comp_A4_350, comp_A1_738, comp_A997_319, comp_A7_411, comp_A4_400, comp_A9992_93, comp_A99994_781, comp_A93_726, comp_A9998_769, comp_A7_415, comp_A9991_972, comp_A993_608, comp_A3_284, comp_A9995_876, comp_A9_859, comp_A9992_129, comp_A3_102, comp_A3_79, comp_A9993_585, comp_A3_124, comp_A91_239, comp_A93_116, comp_A9_811, comp_A3_757, comp_A99991_336, comp_A98_66, comp_A99995_631, comp_A999_732, comp_A9996_244, comp_A995_167, comp_A98_171, comp_A3_981, comp_A9_827, comp_A9992_357, comp_A4_739, comp_A2_876, comp_A99996_412, comp_A9996_202, comp_A9993_525, comp_A7_666, comp_A92_519, comp_A99994_745, comp_A998_448, comp_A9997_490, comp_A9996_448, comp_A997_332, comp_A4_495, comp_A94_29, comp_A7_919, comp_A99997_247, comp_A993_764, comp_A9991_914, comp_A96_609, comp_A9999_832, comp_A99998_189, comp_A996_296, comp_A99999_409, comp_A99994_713, comp_A993_839, comp_A99997_833, comp_A5_327, comp_A2_894, comp_A3_587, comp_A93_629, comp_A999991_302, comp_A99997_824, comp_A9_155, comp_A5_170, comp_A97_991, comp_A995_114, comp_A5_586, comp_A98_162, comp_A991_728, comp_A9996_782, comp_A99992_505, comp_A9995_733, comp_A9991_1016, comp_A9_152, comp_A5_126, comp_A999992_426, comp_A9_784, comp_A999992_487, comp_A92_504, comp_A9994_769, comp_A95_435, comp_A999992_569, comp_A1_652, comp_A991_268, comp_A99997_799, comp_A992_599, comp_A99991_539, comp_A98_147, comp_A7_591, comp_A997_589, comp_A97_124, comp_A996_225, comp_A97_121, comp_A99995_671, comp_A9998_723, comp_A999993_9, comp_A996_92, comp_A996_222, comp_A9999_756, comp_A95_203, comp_A997_838, comp_A5_478, comp_A99997_254, comp_A99991_618, comp_A91_963, comp_A9994_288, comp_A9991_935, comp_A99997_931, comp_A98_151, comp_A4_486, comp_A3_232, comp_A9995_839, comp_A7_592, comp_A3_286, comp_A99999_486, comp_A9991_932, comp_A996_372, comp_A9_156, comp_A7_804, comp_A6_255, comp_A99991_344, comp_A8_757, comp_A993_555, comp_A999994_442, comp_A99992_671, comp_A991_479, comp_A97_610, comp_A999991_570, comp_A9_816, comp_A3_80, comp_A8_822, comp_A998_424, comp_A999993_8, comp_A9992_421, comp_A99999_549, comp_A9993_307, comp_A9996_562, comp_A996_271, comp_A992_400, comp_A94_31, comp_A99_8, comp_A3_54, comp_A2_872, comp_A92_972, comp_A3_272, comp_A999995_1015, comp_A7_605, comp_A9993_295, comp_A991_531, comp_A993_317, comp_A991_869, comp_A94_50, comp_A99994_178, comp_A8_786, comp_A3_407, comp_A6_722, comp_A99999_735, comp_A92_259, comp_A999996_390, comp_A2_901, comp_A992_675, comp_A9_821, comp_A92_503, comp_A8_536, comp_A2_124, comp_A92_250, comp_A95_497, comp_A6_406, comp_A9991_948, comp_A9999_819, comp_A3_535, comp_A998_805, comp_A92_995, comp_A9996_600, comp_A6_606, comp_A996_353, comp_A99994_600, comp_A99991_286, comp_A996_340, comp_A998_414, comp_A996_331, comp_A994_640, comp_A999_714, comp_A3_233, comp_A9_805, comp_A8_540, comp_A99996_575, comp_A993_982, comp_A9993_530, comp_A994_475, comp_A996_332, comp_A4_484, comp_A98_325, comp_A993_659, comp_A2_602, comp_A92_505, comp_A99999_58, comp_A9992_123, comp_A999992_527, comp_A9996_758, comp_A997_428, comp_A3_515, comp_A992_389, comp_A93_513, comp_A99999_558, comp_A9992_429, comp_A993_440, comp_A99996_766, comp_A999991_485, comp_A9991_1009, comp_A99999_594, comp_A993_492, comp_A96_754, comp_A993_321, comp_A999_712, comp_A997_421, comp_A9999_805, comp_A995_343, comp_A9996_570, comp_A5_653, comp_A4_445, comp_A99995_511, comp_A99991_185, comp_A99999_517, comp_A8_334, comp_A9996_737, comp_A9_845, comp_A997_339, comp_A997_243, comp_A993_683, comp_A994_543, comp_A99_13, comp_A2_22, comp_A96_818, comp_A3_350, comp_A992_528, comp_A96_271, comp_A994_365, comp_A999991_372, comp_A99999_168, comp_A95_430, comp_A8_398, comp_A994_484, comp_A999997_1009, comp_A3_415, comp_A97_174, comp_A997_549, comp_A999996_427, comp_A3_381, comp_A997_496, comp_A995_61, comp_A99_15, comp_A99_18, comp_A992_721, comp_A6_474, comp_A95_345, comp_A2_860, comp_A9_853, comp_A93_136, comp_A991_746, comp_A2_320, comp_A97_182, comp_A91_383, comp_A6_485, comp_A99995_471, comp_A93_516, comp_A99992_501, comp_A2_920, comp_A9991_961, comp_A999996_360, comp_A996_350, comp_A991_868, comp_A992_266, comp_A95_312, comp_A96_171, comp_A98_61, comp_A9994_693, comp_A994_378, comp_A99991_182, comp_A8_718, comp_A3_428, comp_A99996_862, comp_A9993_327, comp_A995_537, comp_A9_832, comp_A6_442, comp_A999996_428, comp_A94_58, comp_A997_521, comp_A996_360, comp_A99992_503, comp_A999994_457, comp_A99992_710, comp_A99991_366, comp_A993_286, comp_A999_567, comp_A99996_858, comp_A5_316, comp_A995_299, comp_A991_852, comp_A94_49, comp_A9992_105, comp_A92_247, comp_A98_68, comp_A99995_519, comp_A92_989, comp_A3_285, comp_A94_42, comp_A97_400, comp_A3_209, comp_A8_381, comp_A99_19, comp_A999997_1011, comp_A92_815, comp_A94_33, comp_A9991_937, comp_A998_499, comp_A1_554, comp_A999994_662, comp_A5_562, comp_A9997_669, comp_A997_477, comp_A9991_973, comp_A9999_248, comp_A996_245, comp_A98_1019, comp_A3_112, comp_A994_355, comp_A993_548, comp_A9991_817, comp_A92_246, comp_A3_27, comp_A8_810, comp_A99994_682, comp_A993_612, comp_A9992_99, comp_A9996_610, comp_A997_620, comp_A994_477, comp_A9999_293, comp_A8_404, comp_A996_318, comp_A95_274, comp_A1_601, comp_A92_562, comp_A99997_252, comp_A9996_694, comp_A3_305, comp_A997_334, comp_A999994_507, comp_A99993_647, comp_A992_308, comp_A99992_810, comp_A9993_652, comp_A997_403, comp_A93_651, comp_A999991_306, comp_A991_720, comp_A9992_107, comp_A9_851, comp_A9992_103, comp_A2_869, comp_A997_578, comp_A998_302, comp_A99991_660, comp_A6_644, comp_A2_285, comp_A995_202, comp_A8_818, comp_A999995_1012, comp_A997_956, comp_A999992_388, comp_A93_687, comp_A999995_1008, comp_A996_292, comp_A991_250, comp_A95_354, comp_A9994_711, comp_A9994_295, comp_A5_505, comp_A94_35, comp_A999994_547, comp_A9993_685, comp_A93_718, comp_A9991_956, comp_A993_484, comp_A1_708, comp_A9991_990, comp_A3_283, comp_A998_641, comp_A92_377, comp_A99994_383, comp_A999992_484, comp_A9_160, comp_A997_422, comp_A2_862, comp_A96_180, comp_A99997_843, comp_A9994_704, comp_A98_240, comp_A3_992, comp_A9994_881, comp_A2_827, comp_A999997_1012, comp_A994_549, comp_A97_171, comp_A9993_313, comp_A4_545, comp_A996_200, comp_A3_247, comp_A995_185, comp_A998_559, comp_A9999_767, comp_A99996_551, comp_A6_701, comp_A992_817, comp_A93_115, comp_A9991_962, comp_A99993_596, comp_A93_98, comp_A99994_807, comp_A96_264, comp_A92_500, comp_A9996_693, comp_A99993_630, comp_A99996_513, comp_A997_451, comp_A9992_161, comp_A2_114, comp_A995_493, comp_A99996_188, comp_A3_116, comp_A99996_839, comp_A2_9, comp_A93_544, comp_A3_812, comp_A997_373, comp_A99999_423, comp_A9991_955, comp_A9998_906, comp_A999996_461, comp_A999_585, comp_A5_753, comp_A99993_51, comp_A92_255, comp_A7_856, comp_A9_829, comp_A99995_559, comp_A2_33, comp_A99999_545, comp_A9992_436, comp_A997_666, comp_A94_37, comp_A9991_1011, comp_A99991_408, comp_A996_343, comp_A9999_560, comp_A996_263, comp_A9996_763, comp_A99992_660, comp_A1_642, comp_A9999_419, comp_A7_643, comp_A99992_736, comp_A9_61, comp_A6_394, comp_A99999_406, comp_A3_565, comp_A997_381, comp_A99992_538, comp_A99994_755, comp_A8_484, comp_A99992_655, comp_A991_451, comp_A99995_531, comp_A3_386, comp_A9998_389, comp_A994_390, comp_A97_201, comp_A3_750, comp_A995_34, comp_A994_677, comp_A93_720, comp_A99997_149, comp_A3_588, comp_A98_120, comp_A9_151, comp_A996_244, comp_A9999_786, comp_A99992_744, comp_A97_968, comp_A9993_626, comp_A99998_187, comp_A99994_612, comp_A9991_982, comp_A2_918, comp_A996_304, comp_A99_5, comp_A9991_693, comp_A99_21, comp_A9991_931, comp_A3_103, comp_A998_676, comp_A9_486, comp_A92_528, comp_A7_460, comp_A999994_411, comp_A93_722, comp_A98_153, comp_A996_231, comp_A999_516, comp_A991_373, comp_A9993_658, comp_A999992_474, comp_A999995_1014, comp_A9995_441, comp_A996_327, comp_A1_684, comp_A99999_443, comp_A9996_623, comp_A9_150, comp_A997_713, comp_A9991_965, comp_A999992_432, comp_A999996_726, comp_A993_258, comp_A8_335, comp_A999_656, comp_A991_735, comp_A996_203, comp_A93_546, comp_A99996_508, comp_A99996_263, comp_A9996_431, comp_A96_22, comp_A94_30, comp_A999_711, comp_A9_840, comp_A91_210, comp_A9997_587, comp_A2_713, comp_A999996_685, comp_A2_844, comp_A997_399, comp_A9993_561, comp_A991_391, comp_A6_286, comp_A99992_711, comp_A9991_921, comp_A3_55, comp_A9_157, comp_A8_657, comp_A99994_586, comp_A991_797, comp_A997_394, comp_A96_766, comp_A9993_581, comp_A9998_661, comp_A99993_699, comp_A9996_707, comp_A99997_955, comp_A991_647, comp_A996_185, comp_A999992_536, comp_A93_92, comp_A1_581, comp_A991_486, comp_A993_621, comp_A999992_339, comp_A7_767, comp_A99993_85, comp_A92_574, comp_A3_867, comp_A98_270, comp_A93_119, comp_A992_234, comp_A92_992, comp_A991_644, comp_A3_662, comp_A996_311, comp_A994_457, comp_A9993_539, comp_A99997_946, comp_A997_299, comp_A99992_670, comp_A94_32, comp_A1_741, comp_A994_524, comp_A9997_340, comp_A997_696, comp_A99994_727, comp_A994_644, comp_A996_369, comp_A9991_995, comp_A5_492, comp_A998_230, comp_A93_532, comp_A999_337, comp_A95_388, comp_A3_127, comp_A6_452, comp_A4_332, comp_A999996_581, comp_A8_875, comp_A97_207, comp_A9993_671, comp_A9999_59, comp_A991_777, comp_A9991_699
);

input [9:0] reg_A1;
input [9:0] reg_A2;
input [9:0] reg_A3;
input [9:0] reg_A4;
input [9:0] reg_A5;
input [9:0] reg_A6;
input [9:0] reg_A7;
input [9:0] reg_A8;
input [9:0] reg_A9;
input [9:0] reg_A91;
input [9:0] reg_A92;
input [9:0] reg_A93;
input [9:0] reg_A94;
input [9:0] reg_A95;
input [9:0] reg_A96;
input [9:0] reg_A97;
input [9:0] reg_A98;
input [9:0] reg_A99;
input [9:0] reg_A991;
input [9:0] reg_A992;
input [9:0] reg_A993;
input [9:0] reg_A994;
input [9:0] reg_A995;
input [9:0] reg_A996;
input [9:0] reg_A997;
input [9:0] reg_A998;
input [9:0] reg_A999;
input [9:0] reg_A9991;
input [9:0] reg_A9992;
input [9:0] reg_A9993;
input [9:0] reg_A9994;
input [9:0] reg_A9995;
input [9:0] reg_A9996;
input [9:0] reg_A9997;
input [9:0] reg_A9998;
input [9:0] reg_A9999;
input [9:0] reg_A99991;
input [9:0] reg_A99992;
input [9:0] reg_A99993;
input [9:0] reg_A99994;
input [9:0] reg_A99995;
input [9:0] reg_A99996;
input [9:0] reg_A99997;
input [9:0] reg_A99998;
input [9:0] reg_A99999;
input [9:0] reg_A999991;
input [9:0] reg_A999992;
input [9:0] reg_A999993;
input [9:0] reg_A999994;
input [9:0] reg_A999995;
input [9:0] reg_A999996;
input [9:0] reg_A999997;
output [0:0] comp_A1_649;
output [0:0] comp_A2_29;
output [0:0] comp_A3_322;
output [0:0] comp_A4_504;
output [0:0] comp_A5_495;
output [0:0] comp_A6_624;
output [0:0] comp_A7_593;
output [0:0] comp_A1_220;
output [0:0] comp_A4_472;
output [0:0] comp_A8_701;
output [0:0] comp_A9_178;
output [0:0] comp_A91_362;
output [0:0] comp_A92_263;
output [0:0] comp_A93_529;
output [0:0] comp_A94_40;
output [0:0] comp_A7_795;
output [0:0] comp_A95_118;
output [0:0] comp_A3_541;
output [0:0] comp_A8_90;
output [0:0] comp_A96_11;
output [0:0] comp_A97_193;
output [0:0] comp_A98_202;
output [0:0] comp_A99_14;
output [0:0] comp_A2_830;
output [0:0] comp_A991_288;
output [0:0] comp_A992_452;
output [0:0] comp_A95_373;
output [0:0] comp_A8_777;
output [0:0] comp_A93_537;
output [0:0] comp_A99_11;
output [0:0] comp_A95_383;
output [0:0] comp_A993_454;
output [0:0] comp_A992_774;
output [0:0] comp_A994_302;
output [0:0] comp_A995_87;
output [0:0] comp_A98_143;
output [0:0] comp_A996_348;
output [0:0] comp_A997_750;
output [0:0] comp_A1_884;
output [0:0] comp_A997_360;
output [0:0] comp_A998_765;
output [0:0] comp_A8_726;
output [0:0] comp_A999_643;
output [0:0] comp_A3_526;
output [0:0] comp_A7_455;
output [0:0] comp_A9991_920;
output [0:0] comp_A3_300;
output [0:0] comp_A92_262;
output [0:0] comp_A9992_183;
output [0:0] comp_A991_737;
output [0:0] comp_A97_140;
output [0:0] comp_A9991_923;
output [0:0] comp_A96_873;
output [0:0] comp_A9993_513;
output [0:0] comp_A4_515;
output [0:0] comp_A9994_577;
output [0:0] comp_A94_46;
output [0:0] comp_A7_341;
output [0:0] comp_A3_687;
output [0:0] comp_A9995_483;
output [0:0] comp_A9996_660;
output [0:0] comp_A9997_526;
output [0:0] comp_A9991_943;
output [0:0] comp_A7_561;
output [0:0] comp_A993_276;
output [0:0] comp_A9998_478;
output [0:0] comp_A92_975;
output [0:0] comp_A1_727;
output [0:0] comp_A7_583;
output [0:0] comp_A995_79;
output [0:0] comp_A97_173;
output [0:0] comp_A993_665;
output [0:0] comp_A9999_801;
output [0:0] comp_A3_536;
output [0:0] comp_A999_620;
output [0:0] comp_A994_700;
output [0:0] comp_A99991_242;
output [0:0] comp_A994_712;
output [0:0] comp_A99992_806;
output [0:0] comp_A9997_570;
output [0:0] comp_A99993_119;
output [0:0] comp_A6_670;
output [0:0] comp_A994_338;
output [0:0] comp_A6_635;
output [0:0] comp_A9994_627;
output [0:0] comp_A1_881;
output [0:0] comp_A4_490;
output [0:0] comp_A92_264;
output [0:0] comp_A2_839;
output [0:0] comp_A991_760;
output [0:0] comp_A993_680;
output [0:0] comp_A99994_810;
output [0:0] comp_A98_974;
output [0:0] comp_A4_350;
output [0:0] comp_A1_738;
output [0:0] comp_A997_319;
output [0:0] comp_A7_411;
output [0:0] comp_A4_400;
output [0:0] comp_A9992_93;
output [0:0] comp_A99994_781;
output [0:0] comp_A93_726;
output [0:0] comp_A9998_769;
output [0:0] comp_A7_415;
output [0:0] comp_A9991_972;
output [0:0] comp_A993_608;
output [0:0] comp_A3_284;
output [0:0] comp_A9995_876;
output [0:0] comp_A9_859;
output [0:0] comp_A9992_129;
output [0:0] comp_A3_102;
output [0:0] comp_A3_79;
output [0:0] comp_A9993_585;
output [0:0] comp_A3_124;
output [0:0] comp_A91_239;
output [0:0] comp_A93_116;
output [0:0] comp_A9_811;
output [0:0] comp_A3_757;
output [0:0] comp_A99991_336;
output [0:0] comp_A98_66;
output [0:0] comp_A99995_631;
output [0:0] comp_A999_732;
output [0:0] comp_A9996_244;
output [0:0] comp_A995_167;
output [0:0] comp_A98_171;
output [0:0] comp_A3_981;
output [0:0] comp_A9_827;
output [0:0] comp_A9992_357;
output [0:0] comp_A4_739;
output [0:0] comp_A2_876;
output [0:0] comp_A99996_412;
output [0:0] comp_A9996_202;
output [0:0] comp_A9993_525;
output [0:0] comp_A7_666;
output [0:0] comp_A92_519;
output [0:0] comp_A99994_745;
output [0:0] comp_A998_448;
output [0:0] comp_A9997_490;
output [0:0] comp_A9996_448;
output [0:0] comp_A997_332;
output [0:0] comp_A4_495;
output [0:0] comp_A94_29;
output [0:0] comp_A7_919;
output [0:0] comp_A99997_247;
output [0:0] comp_A993_764;
output [0:0] comp_A9991_914;
output [0:0] comp_A96_609;
output [0:0] comp_A9999_832;
output [0:0] comp_A99998_189;
output [0:0] comp_A996_296;
output [0:0] comp_A99999_409;
output [0:0] comp_A99994_713;
output [0:0] comp_A993_839;
output [0:0] comp_A99997_833;
output [0:0] comp_A5_327;
output [0:0] comp_A2_894;
output [0:0] comp_A3_587;
output [0:0] comp_A93_629;
output [0:0] comp_A999991_302;
output [0:0] comp_A99997_824;
output [0:0] comp_A9_155;
output [0:0] comp_A5_170;
output [0:0] comp_A97_991;
output [0:0] comp_A995_114;
output [0:0] comp_A5_586;
output [0:0] comp_A98_162;
output [0:0] comp_A991_728;
output [0:0] comp_A9996_782;
output [0:0] comp_A99992_505;
output [0:0] comp_A9995_733;
output [0:0] comp_A9991_1016;
output [0:0] comp_A9_152;
output [0:0] comp_A5_126;
output [0:0] comp_A999992_426;
output [0:0] comp_A9_784;
output [0:0] comp_A999992_487;
output [0:0] comp_A92_504;
output [0:0] comp_A9994_769;
output [0:0] comp_A95_435;
output [0:0] comp_A999992_569;
output [0:0] comp_A1_652;
output [0:0] comp_A991_268;
output [0:0] comp_A99997_799;
output [0:0] comp_A992_599;
output [0:0] comp_A99991_539;
output [0:0] comp_A98_147;
output [0:0] comp_A7_591;
output [0:0] comp_A997_589;
output [0:0] comp_A97_124;
output [0:0] comp_A996_225;
output [0:0] comp_A97_121;
output [0:0] comp_A99995_671;
output [0:0] comp_A9998_723;
output [0:0] comp_A999993_9;
output [0:0] comp_A996_92;
output [0:0] comp_A996_222;
output [0:0] comp_A9999_756;
output [0:0] comp_A95_203;
output [0:0] comp_A997_838;
output [0:0] comp_A5_478;
output [0:0] comp_A99997_254;
output [0:0] comp_A99991_618;
output [0:0] comp_A91_963;
output [0:0] comp_A9994_288;
output [0:0] comp_A9991_935;
output [0:0] comp_A99997_931;
output [0:0] comp_A98_151;
output [0:0] comp_A4_486;
output [0:0] comp_A3_232;
output [0:0] comp_A9995_839;
output [0:0] comp_A7_592;
output [0:0] comp_A3_286;
output [0:0] comp_A99999_486;
output [0:0] comp_A9991_932;
output [0:0] comp_A996_372;
output [0:0] comp_A9_156;
output [0:0] comp_A7_804;
output [0:0] comp_A6_255;
output [0:0] comp_A99991_344;
output [0:0] comp_A8_757;
output [0:0] comp_A993_555;
output [0:0] comp_A999994_442;
output [0:0] comp_A99992_671;
output [0:0] comp_A991_479;
output [0:0] comp_A97_610;
output [0:0] comp_A999991_570;
output [0:0] comp_A9_816;
output [0:0] comp_A3_80;
output [0:0] comp_A8_822;
output [0:0] comp_A998_424;
output [0:0] comp_A999993_8;
output [0:0] comp_A9992_421;
output [0:0] comp_A99999_549;
output [0:0] comp_A9993_307;
output [0:0] comp_A9996_562;
output [0:0] comp_A996_271;
output [0:0] comp_A992_400;
output [0:0] comp_A94_31;
output [0:0] comp_A99_8;
output [0:0] comp_A3_54;
output [0:0] comp_A2_872;
output [0:0] comp_A92_972;
output [0:0] comp_A3_272;
output [0:0] comp_A999995_1015;
output [0:0] comp_A7_605;
output [0:0] comp_A9993_295;
output [0:0] comp_A991_531;
output [0:0] comp_A993_317;
output [0:0] comp_A991_869;
output [0:0] comp_A94_50;
output [0:0] comp_A99994_178;
output [0:0] comp_A8_786;
output [0:0] comp_A3_407;
output [0:0] comp_A6_722;
output [0:0] comp_A99999_735;
output [0:0] comp_A92_259;
output [0:0] comp_A999996_390;
output [0:0] comp_A2_901;
output [0:0] comp_A992_675;
output [0:0] comp_A9_821;
output [0:0] comp_A92_503;
output [0:0] comp_A8_536;
output [0:0] comp_A2_124;
output [0:0] comp_A92_250;
output [0:0] comp_A95_497;
output [0:0] comp_A6_406;
output [0:0] comp_A9991_948;
output [0:0] comp_A9999_819;
output [0:0] comp_A3_535;
output [0:0] comp_A998_805;
output [0:0] comp_A92_995;
output [0:0] comp_A9996_600;
output [0:0] comp_A6_606;
output [0:0] comp_A996_353;
output [0:0] comp_A99994_600;
output [0:0] comp_A99991_286;
output [0:0] comp_A996_340;
output [0:0] comp_A998_414;
output [0:0] comp_A996_331;
output [0:0] comp_A994_640;
output [0:0] comp_A999_714;
output [0:0] comp_A3_233;
output [0:0] comp_A9_805;
output [0:0] comp_A8_540;
output [0:0] comp_A99996_575;
output [0:0] comp_A993_982;
output [0:0] comp_A9993_530;
output [0:0] comp_A994_475;
output [0:0] comp_A996_332;
output [0:0] comp_A4_484;
output [0:0] comp_A98_325;
output [0:0] comp_A993_659;
output [0:0] comp_A2_602;
output [0:0] comp_A92_505;
output [0:0] comp_A99999_58;
output [0:0] comp_A9992_123;
output [0:0] comp_A999992_527;
output [0:0] comp_A9996_758;
output [0:0] comp_A997_428;
output [0:0] comp_A3_515;
output [0:0] comp_A992_389;
output [0:0] comp_A93_513;
output [0:0] comp_A99999_558;
output [0:0] comp_A9992_429;
output [0:0] comp_A993_440;
output [0:0] comp_A99996_766;
output [0:0] comp_A999991_485;
output [0:0] comp_A9991_1009;
output [0:0] comp_A99999_594;
output [0:0] comp_A993_492;
output [0:0] comp_A96_754;
output [0:0] comp_A993_321;
output [0:0] comp_A999_712;
output [0:0] comp_A997_421;
output [0:0] comp_A9999_805;
output [0:0] comp_A995_343;
output [0:0] comp_A9996_570;
output [0:0] comp_A5_653;
output [0:0] comp_A4_445;
output [0:0] comp_A99995_511;
output [0:0] comp_A99991_185;
output [0:0] comp_A99999_517;
output [0:0] comp_A8_334;
output [0:0] comp_A9996_737;
output [0:0] comp_A9_845;
output [0:0] comp_A997_339;
output [0:0] comp_A997_243;
output [0:0] comp_A993_683;
output [0:0] comp_A994_543;
output [0:0] comp_A99_13;
output [0:0] comp_A2_22;
output [0:0] comp_A96_818;
output [0:0] comp_A3_350;
output [0:0] comp_A992_528;
output [0:0] comp_A96_271;
output [0:0] comp_A994_365;
output [0:0] comp_A999991_372;
output [0:0] comp_A99999_168;
output [0:0] comp_A95_430;
output [0:0] comp_A8_398;
output [0:0] comp_A994_484;
output [0:0] comp_A999997_1009;
output [0:0] comp_A3_415;
output [0:0] comp_A97_174;
output [0:0] comp_A997_549;
output [0:0] comp_A999996_427;
output [0:0] comp_A3_381;
output [0:0] comp_A997_496;
output [0:0] comp_A995_61;
output [0:0] comp_A99_15;
output [0:0] comp_A99_18;
output [0:0] comp_A992_721;
output [0:0] comp_A6_474;
output [0:0] comp_A95_345;
output [0:0] comp_A2_860;
output [0:0] comp_A9_853;
output [0:0] comp_A93_136;
output [0:0] comp_A991_746;
output [0:0] comp_A2_320;
output [0:0] comp_A97_182;
output [0:0] comp_A91_383;
output [0:0] comp_A6_485;
output [0:0] comp_A99995_471;
output [0:0] comp_A93_516;
output [0:0] comp_A99992_501;
output [0:0] comp_A2_920;
output [0:0] comp_A9991_961;
output [0:0] comp_A999996_360;
output [0:0] comp_A996_350;
output [0:0] comp_A991_868;
output [0:0] comp_A992_266;
output [0:0] comp_A95_312;
output [0:0] comp_A96_171;
output [0:0] comp_A98_61;
output [0:0] comp_A9994_693;
output [0:0] comp_A994_378;
output [0:0] comp_A99991_182;
output [0:0] comp_A8_718;
output [0:0] comp_A3_428;
output [0:0] comp_A99996_862;
output [0:0] comp_A9993_327;
output [0:0] comp_A995_537;
output [0:0] comp_A9_832;
output [0:0] comp_A6_442;
output [0:0] comp_A999996_428;
output [0:0] comp_A94_58;
output [0:0] comp_A997_521;
output [0:0] comp_A996_360;
output [0:0] comp_A99992_503;
output [0:0] comp_A999994_457;
output [0:0] comp_A99992_710;
output [0:0] comp_A99991_366;
output [0:0] comp_A993_286;
output [0:0] comp_A999_567;
output [0:0] comp_A99996_858;
output [0:0] comp_A5_316;
output [0:0] comp_A995_299;
output [0:0] comp_A991_852;
output [0:0] comp_A94_49;
output [0:0] comp_A9992_105;
output [0:0] comp_A92_247;
output [0:0] comp_A98_68;
output [0:0] comp_A99995_519;
output [0:0] comp_A92_989;
output [0:0] comp_A3_285;
output [0:0] comp_A94_42;
output [0:0] comp_A97_400;
output [0:0] comp_A3_209;
output [0:0] comp_A8_381;
output [0:0] comp_A99_19;
output [0:0] comp_A999997_1011;
output [0:0] comp_A92_815;
output [0:0] comp_A94_33;
output [0:0] comp_A9991_937;
output [0:0] comp_A998_499;
output [0:0] comp_A1_554;
output [0:0] comp_A999994_662;
output [0:0] comp_A5_562;
output [0:0] comp_A9997_669;
output [0:0] comp_A997_477;
output [0:0] comp_A9991_973;
output [0:0] comp_A9999_248;
output [0:0] comp_A996_245;
output [0:0] comp_A98_1019;
output [0:0] comp_A3_112;
output [0:0] comp_A994_355;
output [0:0] comp_A993_548;
output [0:0] comp_A9991_817;
output [0:0] comp_A92_246;
output [0:0] comp_A3_27;
output [0:0] comp_A8_810;
output [0:0] comp_A99994_682;
output [0:0] comp_A993_612;
output [0:0] comp_A9992_99;
output [0:0] comp_A9996_610;
output [0:0] comp_A997_620;
output [0:0] comp_A994_477;
output [0:0] comp_A9999_293;
output [0:0] comp_A8_404;
output [0:0] comp_A996_318;
output [0:0] comp_A95_274;
output [0:0] comp_A1_601;
output [0:0] comp_A92_562;
output [0:0] comp_A99997_252;
output [0:0] comp_A9996_694;
output [0:0] comp_A3_305;
output [0:0] comp_A997_334;
output [0:0] comp_A999994_507;
output [0:0] comp_A99993_647;
output [0:0] comp_A992_308;
output [0:0] comp_A99992_810;
output [0:0] comp_A9993_652;
output [0:0] comp_A997_403;
output [0:0] comp_A93_651;
output [0:0] comp_A999991_306;
output [0:0] comp_A991_720;
output [0:0] comp_A9992_107;
output [0:0] comp_A9_851;
output [0:0] comp_A9992_103;
output [0:0] comp_A2_869;
output [0:0] comp_A997_578;
output [0:0] comp_A998_302;
output [0:0] comp_A99991_660;
output [0:0] comp_A6_644;
output [0:0] comp_A2_285;
output [0:0] comp_A995_202;
output [0:0] comp_A8_818;
output [0:0] comp_A999995_1012;
output [0:0] comp_A997_956;
output [0:0] comp_A999992_388;
output [0:0] comp_A93_687;
output [0:0] comp_A999995_1008;
output [0:0] comp_A996_292;
output [0:0] comp_A991_250;
output [0:0] comp_A95_354;
output [0:0] comp_A9994_711;
output [0:0] comp_A9994_295;
output [0:0] comp_A5_505;
output [0:0] comp_A94_35;
output [0:0] comp_A999994_547;
output [0:0] comp_A9993_685;
output [0:0] comp_A93_718;
output [0:0] comp_A9991_956;
output [0:0] comp_A993_484;
output [0:0] comp_A1_708;
output [0:0] comp_A9991_990;
output [0:0] comp_A3_283;
output [0:0] comp_A998_641;
output [0:0] comp_A92_377;
output [0:0] comp_A99994_383;
output [0:0] comp_A999992_484;
output [0:0] comp_A9_160;
output [0:0] comp_A997_422;
output [0:0] comp_A2_862;
output [0:0] comp_A96_180;
output [0:0] comp_A99997_843;
output [0:0] comp_A9994_704;
output [0:0] comp_A98_240;
output [0:0] comp_A3_992;
output [0:0] comp_A9994_881;
output [0:0] comp_A2_827;
output [0:0] comp_A999997_1012;
output [0:0] comp_A994_549;
output [0:0] comp_A97_171;
output [0:0] comp_A9993_313;
output [0:0] comp_A4_545;
output [0:0] comp_A996_200;
output [0:0] comp_A3_247;
output [0:0] comp_A995_185;
output [0:0] comp_A998_559;
output [0:0] comp_A9999_767;
output [0:0] comp_A99996_551;
output [0:0] comp_A6_701;
output [0:0] comp_A992_817;
output [0:0] comp_A93_115;
output [0:0] comp_A9991_962;
output [0:0] comp_A99993_596;
output [0:0] comp_A93_98;
output [0:0] comp_A99994_807;
output [0:0] comp_A96_264;
output [0:0] comp_A92_500;
output [0:0] comp_A9996_693;
output [0:0] comp_A99993_630;
output [0:0] comp_A99996_513;
output [0:0] comp_A997_451;
output [0:0] comp_A9992_161;
output [0:0] comp_A2_114;
output [0:0] comp_A995_493;
output [0:0] comp_A99996_188;
output [0:0] comp_A3_116;
output [0:0] comp_A99996_839;
output [0:0] comp_A2_9;
output [0:0] comp_A93_544;
output [0:0] comp_A3_812;
output [0:0] comp_A997_373;
output [0:0] comp_A99999_423;
output [0:0] comp_A9991_955;
output [0:0] comp_A9998_906;
output [0:0] comp_A999996_461;
output [0:0] comp_A999_585;
output [0:0] comp_A5_753;
output [0:0] comp_A99993_51;
output [0:0] comp_A92_255;
output [0:0] comp_A7_856;
output [0:0] comp_A9_829;
output [0:0] comp_A99995_559;
output [0:0] comp_A2_33;
output [0:0] comp_A99999_545;
output [0:0] comp_A9992_436;
output [0:0] comp_A997_666;
output [0:0] comp_A94_37;
output [0:0] comp_A9991_1011;
output [0:0] comp_A99991_408;
output [0:0] comp_A996_343;
output [0:0] comp_A9999_560;
output [0:0] comp_A996_263;
output [0:0] comp_A9996_763;
output [0:0] comp_A99992_660;
output [0:0] comp_A1_642;
output [0:0] comp_A9999_419;
output [0:0] comp_A7_643;
output [0:0] comp_A99992_736;
output [0:0] comp_A9_61;
output [0:0] comp_A6_394;
output [0:0] comp_A99999_406;
output [0:0] comp_A3_565;
output [0:0] comp_A997_381;
output [0:0] comp_A99992_538;
output [0:0] comp_A99994_755;
output [0:0] comp_A8_484;
output [0:0] comp_A99992_655;
output [0:0] comp_A991_451;
output [0:0] comp_A99995_531;
output [0:0] comp_A3_386;
output [0:0] comp_A9998_389;
output [0:0] comp_A994_390;
output [0:0] comp_A97_201;
output [0:0] comp_A3_750;
output [0:0] comp_A995_34;
output [0:0] comp_A994_677;
output [0:0] comp_A93_720;
output [0:0] comp_A99997_149;
output [0:0] comp_A3_588;
output [0:0] comp_A98_120;
output [0:0] comp_A9_151;
output [0:0] comp_A996_244;
output [0:0] comp_A9999_786;
output [0:0] comp_A99992_744;
output [0:0] comp_A97_968;
output [0:0] comp_A9993_626;
output [0:0] comp_A99998_187;
output [0:0] comp_A99994_612;
output [0:0] comp_A9991_982;
output [0:0] comp_A2_918;
output [0:0] comp_A996_304;
output [0:0] comp_A99_5;
output [0:0] comp_A9991_693;
output [0:0] comp_A99_21;
output [0:0] comp_A9991_931;
output [0:0] comp_A3_103;
output [0:0] comp_A998_676;
output [0:0] comp_A9_486;
output [0:0] comp_A92_528;
output [0:0] comp_A7_460;
output [0:0] comp_A999994_411;
output [0:0] comp_A93_722;
output [0:0] comp_A98_153;
output [0:0] comp_A996_231;
output [0:0] comp_A999_516;
output [0:0] comp_A991_373;
output [0:0] comp_A9993_658;
output [0:0] comp_A999992_474;
output [0:0] comp_A999995_1014;
output [0:0] comp_A9995_441;
output [0:0] comp_A996_327;
output [0:0] comp_A1_684;
output [0:0] comp_A99999_443;
output [0:0] comp_A9996_623;
output [0:0] comp_A9_150;
output [0:0] comp_A997_713;
output [0:0] comp_A9991_965;
output [0:0] comp_A999992_432;
output [0:0] comp_A999996_726;
output [0:0] comp_A993_258;
output [0:0] comp_A8_335;
output [0:0] comp_A999_656;
output [0:0] comp_A991_735;
output [0:0] comp_A996_203;
output [0:0] comp_A93_546;
output [0:0] comp_A99996_508;
output [0:0] comp_A99996_263;
output [0:0] comp_A9996_431;
output [0:0] comp_A96_22;
output [0:0] comp_A94_30;
output [0:0] comp_A999_711;
output [0:0] comp_A9_840;
output [0:0] comp_A91_210;
output [0:0] comp_A9997_587;
output [0:0] comp_A2_713;
output [0:0] comp_A999996_685;
output [0:0] comp_A2_844;
output [0:0] comp_A997_399;
output [0:0] comp_A9993_561;
output [0:0] comp_A991_391;
output [0:0] comp_A6_286;
output [0:0] comp_A99992_711;
output [0:0] comp_A9991_921;
output [0:0] comp_A3_55;
output [0:0] comp_A9_157;
output [0:0] comp_A8_657;
output [0:0] comp_A99994_586;
output [0:0] comp_A991_797;
output [0:0] comp_A997_394;
output [0:0] comp_A96_766;
output [0:0] comp_A9993_581;
output [0:0] comp_A9998_661;
output [0:0] comp_A99993_699;
output [0:0] comp_A9996_707;
output [0:0] comp_A99997_955;
output [0:0] comp_A991_647;
output [0:0] comp_A996_185;
output [0:0] comp_A999992_536;
output [0:0] comp_A93_92;
output [0:0] comp_A1_581;
output [0:0] comp_A991_486;
output [0:0] comp_A993_621;
output [0:0] comp_A999992_339;
output [0:0] comp_A7_767;
output [0:0] comp_A99993_85;
output [0:0] comp_A92_574;
output [0:0] comp_A3_867;
output [0:0] comp_A98_270;
output [0:0] comp_A93_119;
output [0:0] comp_A992_234;
output [0:0] comp_A92_992;
output [0:0] comp_A991_644;
output [0:0] comp_A3_662;
output [0:0] comp_A996_311;
output [0:0] comp_A994_457;
output [0:0] comp_A9993_539;
output [0:0] comp_A99997_946;
output [0:0] comp_A997_299;
output [0:0] comp_A99992_670;
output [0:0] comp_A94_32;
output [0:0] comp_A1_741;
output [0:0] comp_A994_524;
output [0:0] comp_A9997_340;
output [0:0] comp_A997_696;
output [0:0] comp_A99994_727;
output [0:0] comp_A994_644;
output [0:0] comp_A996_369;
output [0:0] comp_A9991_995;
output [0:0] comp_A5_492;
output [0:0] comp_A998_230;
output [0:0] comp_A93_532;
output [0:0] comp_A999_337;
output [0:0] comp_A95_388;
output [0:0] comp_A3_127;
output [0:0] comp_A6_452;
output [0:0] comp_A4_332;
output [0:0] comp_A999996_581;
output [0:0] comp_A8_875;
output [0:0] comp_A97_207;
output [0:0] comp_A9993_671;
output [0:0] comp_A9999_59;
output [0:0] comp_A991_777;
output [0:0] comp_A9991_699;

wire [9:0] const_649_10;
assign const_649_10 = 10'b1010001001;
wire [9:0] const_29_10;
assign const_29_10 = 10'b0000011101;
wire [9:0] const_322_10;
assign const_322_10 = 10'b0101000010;
wire [9:0] const_504_10;
assign const_504_10 = 10'b0111111000;
wire [9:0] const_495_10;
assign const_495_10 = 10'b0111101111;
wire [9:0] const_624_10;
assign const_624_10 = 10'b1001110000;
wire [9:0] const_593_10;
assign const_593_10 = 10'b1001010001;
wire [9:0] const_220_10;
assign const_220_10 = 10'b0011011100;
wire [9:0] const_472_10;
assign const_472_10 = 10'b0111011000;
wire [9:0] const_701_10;
assign const_701_10 = 10'b1010111101;
wire [9:0] const_178_10;
assign const_178_10 = 10'b0010110010;
wire [9:0] const_362_10;
assign const_362_10 = 10'b0101101010;
wire [9:0] const_263_10;
assign const_263_10 = 10'b0100000111;
wire [9:0] const_529_10;
assign const_529_10 = 10'b1000010001;
wire [9:0] const_40_10;
assign const_40_10 = 10'b0000101000;
wire [9:0] const_795_10;
assign const_795_10 = 10'b1100011011;
wire [9:0] const_118_10;
assign const_118_10 = 10'b0001110110;
wire [9:0] const_541_10;
assign const_541_10 = 10'b1000011101;
wire [9:0] const_90_10;
assign const_90_10 = 10'b0001011010;
wire [9:0] const_11_10;
assign const_11_10 = 10'b0000001011;
wire [9:0] const_193_10;
assign const_193_10 = 10'b0011000001;
wire [9:0] const_202_10;
assign const_202_10 = 10'b0011001010;
wire [9:0] const_14_10;
assign const_14_10 = 10'b0000001110;
wire [9:0] const_830_10;
assign const_830_10 = 10'b1100111110;
wire [9:0] const_288_10;
assign const_288_10 = 10'b0100100000;
wire [9:0] const_452_10;
assign const_452_10 = 10'b0111000100;
wire [9:0] const_373_10;
assign const_373_10 = 10'b0101110101;
wire [9:0] const_777_10;
assign const_777_10 = 10'b1100001001;
wire [9:0] const_537_10;
assign const_537_10 = 10'b1000011001;
wire [9:0] const_383_10;
assign const_383_10 = 10'b0101111111;
wire [9:0] const_454_10;
assign const_454_10 = 10'b0111000110;
wire [9:0] const_774_10;
assign const_774_10 = 10'b1100000110;
wire [9:0] const_302_10;
assign const_302_10 = 10'b0100101110;
wire [9:0] const_87_10;
assign const_87_10 = 10'b0001010111;
wire [9:0] const_143_10;
assign const_143_10 = 10'b0010001111;
wire [9:0] const_348_10;
assign const_348_10 = 10'b0101011100;
wire [9:0] const_750_10;
assign const_750_10 = 10'b1011101110;
wire [9:0] const_884_10;
assign const_884_10 = 10'b1101110100;
wire [9:0] const_360_10;
assign const_360_10 = 10'b0101101000;
wire [9:0] const_765_10;
assign const_765_10 = 10'b1011111101;
wire [9:0] const_726_10;
assign const_726_10 = 10'b1011010110;
wire [9:0] const_643_10;
assign const_643_10 = 10'b1010000011;
wire [9:0] const_526_10;
assign const_526_10 = 10'b1000001110;
wire [9:0] const_455_10;
assign const_455_10 = 10'b0111000111;
wire [9:0] const_920_10;
assign const_920_10 = 10'b1110011000;
wire [9:0] const_300_10;
assign const_300_10 = 10'b0100101100;
wire [9:0] const_262_10;
assign const_262_10 = 10'b0100000110;
wire [9:0] const_183_10;
assign const_183_10 = 10'b0010110111;
wire [9:0] const_737_10;
assign const_737_10 = 10'b1011100001;
wire [9:0] const_140_10;
assign const_140_10 = 10'b0010001100;
wire [9:0] const_923_10;
assign const_923_10 = 10'b1110011011;
wire [9:0] const_873_10;
assign const_873_10 = 10'b1101101001;
wire [9:0] const_513_10;
assign const_513_10 = 10'b1000000001;
wire [9:0] const_515_10;
assign const_515_10 = 10'b1000000011;
wire [9:0] const_577_10;
assign const_577_10 = 10'b1001000001;
wire [9:0] const_46_10;
assign const_46_10 = 10'b0000101110;
wire [9:0] const_341_10;
assign const_341_10 = 10'b0101010101;
wire [9:0] const_687_10;
assign const_687_10 = 10'b1010101111;
wire [9:0] const_483_10;
assign const_483_10 = 10'b0111100011;
wire [9:0] const_660_10;
assign const_660_10 = 10'b1010010100;
wire [9:0] const_943_10;
assign const_943_10 = 10'b1110101111;
wire [9:0] const_561_10;
assign const_561_10 = 10'b1000110001;
wire [9:0] const_276_10;
assign const_276_10 = 10'b0100010100;
wire [9:0] const_478_10;
assign const_478_10 = 10'b0111011110;
wire [9:0] const_975_10;
assign const_975_10 = 10'b1111001111;
wire [9:0] const_727_10;
assign const_727_10 = 10'b1011010111;
wire [9:0] const_583_10;
assign const_583_10 = 10'b1001000111;
wire [9:0] const_79_10;
assign const_79_10 = 10'b0001001111;
wire [9:0] const_173_10;
assign const_173_10 = 10'b0010101101;
wire [9:0] const_665_10;
assign const_665_10 = 10'b1010011001;
wire [9:0] const_801_10;
assign const_801_10 = 10'b1100100001;
wire [9:0] const_536_10;
assign const_536_10 = 10'b1000011000;
wire [9:0] const_620_10;
assign const_620_10 = 10'b1001101100;
wire [9:0] const_700_10;
assign const_700_10 = 10'b1010111100;
wire [9:0] const_242_10;
assign const_242_10 = 10'b0011110010;
wire [9:0] const_712_10;
assign const_712_10 = 10'b1011001000;
wire [9:0] const_806_10;
assign const_806_10 = 10'b1100100110;
wire [9:0] const_570_10;
assign const_570_10 = 10'b1000111010;
wire [9:0] const_119_10;
assign const_119_10 = 10'b0001110111;
wire [9:0] const_670_10;
assign const_670_10 = 10'b1010011110;
wire [9:0] const_338_10;
assign const_338_10 = 10'b0101010010;
wire [9:0] const_635_10;
assign const_635_10 = 10'b1001111011;
wire [9:0] const_627_10;
assign const_627_10 = 10'b1001110011;
wire [9:0] const_881_10;
assign const_881_10 = 10'b1101110001;
wire [9:0] const_490_10;
assign const_490_10 = 10'b0111101010;
wire [9:0] const_264_10;
assign const_264_10 = 10'b0100001000;
wire [9:0] const_839_10;
assign const_839_10 = 10'b1101000111;
wire [9:0] const_760_10;
assign const_760_10 = 10'b1011111000;
wire [9:0] const_680_10;
assign const_680_10 = 10'b1010101000;
wire [9:0] const_810_10;
assign const_810_10 = 10'b1100101010;
wire [9:0] const_974_10;
assign const_974_10 = 10'b1111001110;
wire [9:0] const_350_10;
assign const_350_10 = 10'b0101011110;
wire [9:0] const_738_10;
assign const_738_10 = 10'b1011100010;
wire [9:0] const_319_10;
assign const_319_10 = 10'b0100111111;
wire [9:0] const_411_10;
assign const_411_10 = 10'b0110011011;
wire [9:0] const_400_10;
assign const_400_10 = 10'b0110010000;
wire [9:0] const_93_10;
assign const_93_10 = 10'b0001011101;
wire [9:0] const_781_10;
assign const_781_10 = 10'b1100001101;
wire [9:0] const_769_10;
assign const_769_10 = 10'b1100000001;
wire [9:0] const_415_10;
assign const_415_10 = 10'b0110011111;
wire [9:0] const_972_10;
assign const_972_10 = 10'b1111001100;
wire [9:0] const_608_10;
assign const_608_10 = 10'b1001100000;
wire [9:0] const_284_10;
assign const_284_10 = 10'b0100011100;
wire [9:0] const_876_10;
assign const_876_10 = 10'b1101101100;
wire [9:0] const_859_10;
assign const_859_10 = 10'b1101011011;
wire [9:0] const_129_10;
assign const_129_10 = 10'b0010000001;
wire [9:0] const_102_10;
assign const_102_10 = 10'b0001100110;
wire [9:0] const_585_10;
assign const_585_10 = 10'b1001001001;
wire [9:0] const_124_10;
assign const_124_10 = 10'b0001111100;
wire [9:0] const_239_10;
assign const_239_10 = 10'b0011101111;
wire [9:0] const_116_10;
assign const_116_10 = 10'b0001110100;
wire [9:0] const_811_10;
assign const_811_10 = 10'b1100101011;
wire [9:0] const_757_10;
assign const_757_10 = 10'b1011110101;
wire [9:0] const_336_10;
assign const_336_10 = 10'b0101010000;
wire [9:0] const_66_10;
assign const_66_10 = 10'b0001000010;
wire [9:0] const_631_10;
assign const_631_10 = 10'b1001110111;
wire [9:0] const_732_10;
assign const_732_10 = 10'b1011011100;
wire [9:0] const_244_10;
assign const_244_10 = 10'b0011110100;
wire [9:0] const_167_10;
assign const_167_10 = 10'b0010100111;
wire [9:0] const_171_10;
assign const_171_10 = 10'b0010101011;
wire [9:0] const_981_10;
assign const_981_10 = 10'b1111010101;
wire [9:0] const_827_10;
assign const_827_10 = 10'b1100111011;
wire [9:0] const_357_10;
assign const_357_10 = 10'b0101100101;
wire [9:0] const_739_10;
assign const_739_10 = 10'b1011100011;
wire [9:0] const_412_10;
assign const_412_10 = 10'b0110011100;
wire [9:0] const_525_10;
assign const_525_10 = 10'b1000001101;
wire [9:0] const_666_10;
assign const_666_10 = 10'b1010011010;
wire [9:0] const_519_10;
assign const_519_10 = 10'b1000000111;
wire [9:0] const_745_10;
assign const_745_10 = 10'b1011101001;
wire [9:0] const_448_10;
assign const_448_10 = 10'b0111000000;
wire [9:0] const_332_10;
assign const_332_10 = 10'b0101001100;
wire [9:0] const_919_10;
assign const_919_10 = 10'b1110010111;
wire [9:0] const_247_10;
assign const_247_10 = 10'b0011110111;
wire [9:0] const_764_10;
assign const_764_10 = 10'b1011111100;
wire [9:0] const_914_10;
assign const_914_10 = 10'b1110010010;
wire [9:0] const_609_10;
assign const_609_10 = 10'b1001100001;
wire [9:0] const_832_10;
assign const_832_10 = 10'b1101000000;
wire [9:0] const_189_10;
assign const_189_10 = 10'b0010111101;
wire [9:0] const_296_10;
assign const_296_10 = 10'b0100101000;
wire [9:0] const_409_10;
assign const_409_10 = 10'b0110011001;
wire [9:0] const_713_10;
assign const_713_10 = 10'b1011001001;
wire [9:0] const_833_10;
assign const_833_10 = 10'b1101000001;
wire [9:0] const_327_10;
assign const_327_10 = 10'b0101000111;
wire [9:0] const_894_10;
assign const_894_10 = 10'b1101111110;
wire [9:0] const_587_10;
assign const_587_10 = 10'b1001001011;
wire [9:0] const_629_10;
assign const_629_10 = 10'b1001110101;
wire [9:0] const_824_10;
assign const_824_10 = 10'b1100111000;
wire [9:0] const_155_10;
assign const_155_10 = 10'b0010011011;
wire [9:0] const_170_10;
assign const_170_10 = 10'b0010101010;
wire [9:0] const_991_10;
assign const_991_10 = 10'b1111011111;
wire [9:0] const_114_10;
assign const_114_10 = 10'b0001110010;
wire [9:0] const_586_10;
assign const_586_10 = 10'b1001001010;
wire [9:0] const_162_10;
assign const_162_10 = 10'b0010100010;
wire [9:0] const_728_10;
assign const_728_10 = 10'b1011011000;
wire [9:0] const_782_10;
assign const_782_10 = 10'b1100001110;
wire [9:0] const_505_10;
assign const_505_10 = 10'b0111111001;
wire [9:0] const_733_10;
assign const_733_10 = 10'b1011011101;
wire [9:0] const_1016_10;
assign const_1016_10 = 10'b1111111000;
wire [9:0] const_152_10;
assign const_152_10 = 10'b0010011000;
wire [9:0] const_126_10;
assign const_126_10 = 10'b0001111110;
wire [9:0] const_426_10;
assign const_426_10 = 10'b0110101010;
wire [9:0] const_784_10;
assign const_784_10 = 10'b1100010000;
wire [9:0] const_487_10;
assign const_487_10 = 10'b0111100111;
wire [9:0] const_435_10;
assign const_435_10 = 10'b0110110011;
wire [9:0] const_569_10;
assign const_569_10 = 10'b1000111001;
wire [9:0] const_652_10;
assign const_652_10 = 10'b1010001100;
wire [9:0] const_268_10;
assign const_268_10 = 10'b0100001100;
wire [9:0] const_799_10;
assign const_799_10 = 10'b1100011111;
wire [9:0] const_599_10;
assign const_599_10 = 10'b1001010111;
wire [9:0] const_539_10;
assign const_539_10 = 10'b1000011011;
wire [9:0] const_147_10;
assign const_147_10 = 10'b0010010011;
wire [9:0] const_591_10;
assign const_591_10 = 10'b1001001111;
wire [9:0] const_589_10;
assign const_589_10 = 10'b1001001101;
wire [9:0] const_225_10;
assign const_225_10 = 10'b0011100001;
wire [9:0] const_121_10;
assign const_121_10 = 10'b0001111001;
wire [9:0] const_671_10;
assign const_671_10 = 10'b1010011111;
wire [9:0] const_723_10;
assign const_723_10 = 10'b1011010011;
wire [9:0] const_9_10;
assign const_9_10 = 10'b0000001001;
wire [9:0] const_92_10;
assign const_92_10 = 10'b0001011100;
wire [9:0] const_222_10;
assign const_222_10 = 10'b0011011110;
wire [9:0] const_756_10;
assign const_756_10 = 10'b1011110100;
wire [9:0] const_203_10;
assign const_203_10 = 10'b0011001011;
wire [9:0] const_838_10;
assign const_838_10 = 10'b1101000110;
wire [9:0] const_254_10;
assign const_254_10 = 10'b0011111110;
wire [9:0] const_618_10;
assign const_618_10 = 10'b1001101010;
wire [9:0] const_963_10;
assign const_963_10 = 10'b1111000011;
wire [9:0] const_935_10;
assign const_935_10 = 10'b1110100111;
wire [9:0] const_931_10;
assign const_931_10 = 10'b1110100011;
wire [9:0] const_151_10;
assign const_151_10 = 10'b0010010111;
wire [9:0] const_486_10;
assign const_486_10 = 10'b0111100110;
wire [9:0] const_232_10;
assign const_232_10 = 10'b0011101000;
wire [9:0] const_592_10;
assign const_592_10 = 10'b1001010000;
wire [9:0] const_286_10;
assign const_286_10 = 10'b0100011110;
wire [9:0] const_932_10;
assign const_932_10 = 10'b1110100100;
wire [9:0] const_372_10;
assign const_372_10 = 10'b0101110100;
wire [9:0] const_156_10;
assign const_156_10 = 10'b0010011100;
wire [9:0] const_804_10;
assign const_804_10 = 10'b1100100100;
wire [9:0] const_255_10;
assign const_255_10 = 10'b0011111111;
wire [9:0] const_344_10;
assign const_344_10 = 10'b0101011000;
wire [9:0] const_555_10;
assign const_555_10 = 10'b1000101011;
wire [9:0] const_442_10;
assign const_442_10 = 10'b0110111010;
wire [9:0] const_479_10;
assign const_479_10 = 10'b0111011111;
wire [9:0] const_610_10;
assign const_610_10 = 10'b1001100010;
wire [9:0] const_816_10;
assign const_816_10 = 10'b1100110000;
wire [9:0] const_80_10;
assign const_80_10 = 10'b0001010000;
wire [9:0] const_822_10;
assign const_822_10 = 10'b1100110110;
wire [9:0] const_424_10;
assign const_424_10 = 10'b0110101000;
wire [9:0] const_8_10;
assign const_8_10 = 10'b0000001000;
wire [9:0] const_421_10;
assign const_421_10 = 10'b0110100101;
wire [9:0] const_549_10;
assign const_549_10 = 10'b1000100101;
wire [9:0] const_307_10;
assign const_307_10 = 10'b0100110011;
wire [9:0] const_562_10;
assign const_562_10 = 10'b1000110010;
wire [9:0] const_271_10;
assign const_271_10 = 10'b0100001111;
wire [9:0] const_31_10;
assign const_31_10 = 10'b0000011111;
wire [9:0] const_54_10;
assign const_54_10 = 10'b0000110110;
wire [9:0] const_872_10;
assign const_872_10 = 10'b1101101000;
wire [9:0] const_272_10;
assign const_272_10 = 10'b0100010000;
wire [9:0] const_1015_10;
assign const_1015_10 = 10'b1111110111;
wire [9:0] const_605_10;
assign const_605_10 = 10'b1001011101;
wire [9:0] const_295_10;
assign const_295_10 = 10'b0100100111;
wire [9:0] const_531_10;
assign const_531_10 = 10'b1000010011;
wire [9:0] const_317_10;
assign const_317_10 = 10'b0100111101;
wire [9:0] const_869_10;
assign const_869_10 = 10'b1101100101;
wire [9:0] const_50_10;
assign const_50_10 = 10'b0000110010;
wire [9:0] const_786_10;
assign const_786_10 = 10'b1100010010;
wire [9:0] const_407_10;
assign const_407_10 = 10'b0110010111;
wire [9:0] const_722_10;
assign const_722_10 = 10'b1011010010;
wire [9:0] const_735_10;
assign const_735_10 = 10'b1011011111;
wire [9:0] const_259_10;
assign const_259_10 = 10'b0100000011;
wire [9:0] const_390_10;
assign const_390_10 = 10'b0110000110;
wire [9:0] const_901_10;
assign const_901_10 = 10'b1110000101;
wire [9:0] const_675_10;
assign const_675_10 = 10'b1010100011;
wire [9:0] const_821_10;
assign const_821_10 = 10'b1100110101;
wire [9:0] const_503_10;
assign const_503_10 = 10'b0111110111;
wire [9:0] const_250_10;
assign const_250_10 = 10'b0011111010;
wire [9:0] const_497_10;
assign const_497_10 = 10'b0111110001;
wire [9:0] const_406_10;
assign const_406_10 = 10'b0110010110;
wire [9:0] const_948_10;
assign const_948_10 = 10'b1110110100;
wire [9:0] const_819_10;
assign const_819_10 = 10'b1100110011;
wire [9:0] const_535_10;
assign const_535_10 = 10'b1000010111;
wire [9:0] const_805_10;
assign const_805_10 = 10'b1100100101;
wire [9:0] const_995_10;
assign const_995_10 = 10'b1111100011;
wire [9:0] const_600_10;
assign const_600_10 = 10'b1001011000;
wire [9:0] const_606_10;
assign const_606_10 = 10'b1001011110;
wire [9:0] const_353_10;
assign const_353_10 = 10'b0101100001;
wire [9:0] const_340_10;
assign const_340_10 = 10'b0101010100;
wire [9:0] const_414_10;
assign const_414_10 = 10'b0110011110;
wire [9:0] const_331_10;
assign const_331_10 = 10'b0101001011;
wire [9:0] const_640_10;
assign const_640_10 = 10'b1010000000;
wire [9:0] const_714_10;
assign const_714_10 = 10'b1011001010;
wire [9:0] const_233_10;
assign const_233_10 = 10'b0011101001;
wire [9:0] const_540_10;
assign const_540_10 = 10'b1000011100;
wire [9:0] const_575_10;
assign const_575_10 = 10'b1000111111;
wire [9:0] const_982_10;
assign const_982_10 = 10'b1111010110;
wire [9:0] const_530_10;
assign const_530_10 = 10'b1000010010;
wire [9:0] const_475_10;
assign const_475_10 = 10'b0111011011;
wire [9:0] const_484_10;
assign const_484_10 = 10'b0111100100;
wire [9:0] const_325_10;
assign const_325_10 = 10'b0101000101;
wire [9:0] const_659_10;
assign const_659_10 = 10'b1010010011;
wire [9:0] const_602_10;
assign const_602_10 = 10'b1001011010;
wire [9:0] const_58_10;
assign const_58_10 = 10'b0000111010;
wire [9:0] const_123_10;
assign const_123_10 = 10'b0001111011;
wire [9:0] const_527_10;
assign const_527_10 = 10'b1000001111;
wire [9:0] const_758_10;
assign const_758_10 = 10'b1011110110;
wire [9:0] const_428_10;
assign const_428_10 = 10'b0110101100;
wire [9:0] const_389_10;
assign const_389_10 = 10'b0110000101;
wire [9:0] const_558_10;
assign const_558_10 = 10'b1000101110;
wire [9:0] const_429_10;
assign const_429_10 = 10'b0110101101;
wire [9:0] const_440_10;
assign const_440_10 = 10'b0110111000;
wire [9:0] const_766_10;
assign const_766_10 = 10'b1011111110;
wire [9:0] const_485_10;
assign const_485_10 = 10'b0111100101;
wire [9:0] const_1009_10;
assign const_1009_10 = 10'b1111110001;
wire [9:0] const_594_10;
assign const_594_10 = 10'b1001010010;
wire [9:0] const_492_10;
assign const_492_10 = 10'b0111101100;
wire [9:0] const_754_10;
assign const_754_10 = 10'b1011110010;
wire [9:0] const_321_10;
assign const_321_10 = 10'b0101000001;
wire [9:0] const_343_10;
assign const_343_10 = 10'b0101010111;
wire [9:0] const_653_10;
assign const_653_10 = 10'b1010001101;
wire [9:0] const_445_10;
assign const_445_10 = 10'b0110111101;
wire [9:0] const_511_10;
assign const_511_10 = 10'b0111111111;
wire [9:0] const_185_10;
assign const_185_10 = 10'b0010111001;
wire [9:0] const_517_10;
assign const_517_10 = 10'b1000000101;
wire [9:0] const_334_10;
assign const_334_10 = 10'b0101001110;
wire [9:0] const_845_10;
assign const_845_10 = 10'b1101001101;
wire [9:0] const_339_10;
assign const_339_10 = 10'b0101010011;
wire [9:0] const_243_10;
assign const_243_10 = 10'b0011110011;
wire [9:0] const_683_10;
assign const_683_10 = 10'b1010101011;
wire [9:0] const_543_10;
assign const_543_10 = 10'b1000011111;
wire [9:0] const_13_10;
assign const_13_10 = 10'b0000001101;
wire [9:0] const_22_10;
assign const_22_10 = 10'b0000010110;
wire [9:0] const_818_10;
assign const_818_10 = 10'b1100110010;
wire [9:0] const_528_10;
assign const_528_10 = 10'b1000010000;
wire [9:0] const_365_10;
assign const_365_10 = 10'b0101101101;
wire [9:0] const_168_10;
assign const_168_10 = 10'b0010101000;
wire [9:0] const_430_10;
assign const_430_10 = 10'b0110101110;
wire [9:0] const_398_10;
assign const_398_10 = 10'b0110001110;
wire [9:0] const_174_10;
assign const_174_10 = 10'b0010101110;
wire [9:0] const_427_10;
assign const_427_10 = 10'b0110101011;
wire [9:0] const_381_10;
assign const_381_10 = 10'b0101111101;
wire [9:0] const_496_10;
assign const_496_10 = 10'b0111110000;
wire [9:0] const_61_10;
assign const_61_10 = 10'b0000111101;
wire [9:0] const_15_10;
assign const_15_10 = 10'b0000001111;
wire [9:0] const_18_10;
assign const_18_10 = 10'b0000010010;
wire [9:0] const_721_10;
assign const_721_10 = 10'b1011010001;
wire [9:0] const_474_10;
assign const_474_10 = 10'b0111011010;
wire [9:0] const_345_10;
assign const_345_10 = 10'b0101011001;
wire [9:0] const_860_10;
assign const_860_10 = 10'b1101011100;
wire [9:0] const_853_10;
assign const_853_10 = 10'b1101010101;
wire [9:0] const_136_10;
assign const_136_10 = 10'b0010001000;
wire [9:0] const_746_10;
assign const_746_10 = 10'b1011101010;
wire [9:0] const_320_10;
assign const_320_10 = 10'b0101000000;
wire [9:0] const_182_10;
assign const_182_10 = 10'b0010110110;
wire [9:0] const_471_10;
assign const_471_10 = 10'b0111010111;
wire [9:0] const_516_10;
assign const_516_10 = 10'b1000000100;
wire [9:0] const_501_10;
assign const_501_10 = 10'b0111110101;
wire [9:0] const_961_10;
assign const_961_10 = 10'b1111000001;
wire [9:0] const_868_10;
assign const_868_10 = 10'b1101100100;
wire [9:0] const_266_10;
assign const_266_10 = 10'b0100001010;
wire [9:0] const_312_10;
assign const_312_10 = 10'b0100111000;
wire [9:0] const_693_10;
assign const_693_10 = 10'b1010110101;
wire [9:0] const_378_10;
assign const_378_10 = 10'b0101111010;
wire [9:0] const_718_10;
assign const_718_10 = 10'b1011001110;
wire [9:0] const_862_10;
assign const_862_10 = 10'b1101011110;
wire [9:0] const_521_10;
assign const_521_10 = 10'b1000001001;
wire [9:0] const_457_10;
assign const_457_10 = 10'b0111001001;
wire [9:0] const_710_10;
assign const_710_10 = 10'b1011000110;
wire [9:0] const_366_10;
assign const_366_10 = 10'b0101101110;
wire [9:0] const_567_10;
assign const_567_10 = 10'b1000110111;
wire [9:0] const_858_10;
assign const_858_10 = 10'b1101011010;
wire [9:0] const_316_10;
assign const_316_10 = 10'b0100111100;
wire [9:0] const_299_10;
assign const_299_10 = 10'b0100101011;
wire [9:0] const_852_10;
assign const_852_10 = 10'b1101010100;
wire [9:0] const_49_10;
assign const_49_10 = 10'b0000110001;
wire [9:0] const_105_10;
assign const_105_10 = 10'b0001101001;
wire [9:0] const_68_10;
assign const_68_10 = 10'b0001000100;
wire [9:0] const_989_10;
assign const_989_10 = 10'b1111011101;
wire [9:0] const_285_10;
assign const_285_10 = 10'b0100011101;
wire [9:0] const_42_10;
assign const_42_10 = 10'b0000101010;
wire [9:0] const_209_10;
assign const_209_10 = 10'b0011010001;
wire [9:0] const_19_10;
assign const_19_10 = 10'b0000010011;
wire [9:0] const_1011_10;
assign const_1011_10 = 10'b1111110011;
wire [9:0] const_815_10;
assign const_815_10 = 10'b1100101111;
wire [9:0] const_33_10;
assign const_33_10 = 10'b0000100001;
wire [9:0] const_937_10;
assign const_937_10 = 10'b1110101001;
wire [9:0] const_499_10;
assign const_499_10 = 10'b0111110011;
wire [9:0] const_554_10;
assign const_554_10 = 10'b1000101010;
wire [9:0] const_662_10;
assign const_662_10 = 10'b1010010110;
wire [9:0] const_669_10;
assign const_669_10 = 10'b1010011101;
wire [9:0] const_477_10;
assign const_477_10 = 10'b0111011101;
wire [9:0] const_973_10;
assign const_973_10 = 10'b1111001101;
wire [9:0] const_248_10;
assign const_248_10 = 10'b0011111000;
wire [9:0] const_245_10;
assign const_245_10 = 10'b0011110101;
wire [9:0] const_1019_10;
assign const_1019_10 = 10'b1111111011;
wire [9:0] const_112_10;
assign const_112_10 = 10'b0001110000;
wire [9:0] const_355_10;
assign const_355_10 = 10'b0101100011;
wire [9:0] const_548_10;
assign const_548_10 = 10'b1000100100;
wire [9:0] const_817_10;
assign const_817_10 = 10'b1100110001;
wire [9:0] const_246_10;
assign const_246_10 = 10'b0011110110;
wire [9:0] const_27_10;
assign const_27_10 = 10'b0000011011;
wire [9:0] const_682_10;
assign const_682_10 = 10'b1010101010;
wire [9:0] const_612_10;
assign const_612_10 = 10'b1001100100;
wire [9:0] const_99_10;
assign const_99_10 = 10'b0001100011;
wire [9:0] const_293_10;
assign const_293_10 = 10'b0100100101;
wire [9:0] const_404_10;
assign const_404_10 = 10'b0110010100;
wire [9:0] const_318_10;
assign const_318_10 = 10'b0100111110;
wire [9:0] const_274_10;
assign const_274_10 = 10'b0100010010;
wire [9:0] const_601_10;
assign const_601_10 = 10'b1001011001;
wire [9:0] const_252_10;
assign const_252_10 = 10'b0011111100;
wire [9:0] const_694_10;
assign const_694_10 = 10'b1010110110;
wire [9:0] const_305_10;
assign const_305_10 = 10'b0100110001;
wire [9:0] const_507_10;
assign const_507_10 = 10'b0111111011;
wire [9:0] const_647_10;
assign const_647_10 = 10'b1010000111;
wire [9:0] const_308_10;
assign const_308_10 = 10'b0100110100;
wire [9:0] const_403_10;
assign const_403_10 = 10'b0110010011;
wire [9:0] const_651_10;
assign const_651_10 = 10'b1010001011;
wire [9:0] const_306_10;
assign const_306_10 = 10'b0100110010;
wire [9:0] const_720_10;
assign const_720_10 = 10'b1011010000;
wire [9:0] const_107_10;
assign const_107_10 = 10'b0001101011;
wire [9:0] const_851_10;
assign const_851_10 = 10'b1101010011;
wire [9:0] const_103_10;
assign const_103_10 = 10'b0001100111;
wire [9:0] const_578_10;
assign const_578_10 = 10'b1001000010;
wire [9:0] const_644_10;
assign const_644_10 = 10'b1010000100;
wire [9:0] const_1012_10;
assign const_1012_10 = 10'b1111110100;
wire [9:0] const_956_10;
assign const_956_10 = 10'b1110111100;
wire [9:0] const_388_10;
assign const_388_10 = 10'b0110000100;
wire [9:0] const_1008_10;
assign const_1008_10 = 10'b1111110000;
wire [9:0] const_292_10;
assign const_292_10 = 10'b0100100100;
wire [9:0] const_354_10;
assign const_354_10 = 10'b0101100010;
wire [9:0] const_711_10;
assign const_711_10 = 10'b1011000111;
wire [9:0] const_35_10;
assign const_35_10 = 10'b0000100011;
wire [9:0] const_547_10;
assign const_547_10 = 10'b1000100011;
wire [9:0] const_685_10;
assign const_685_10 = 10'b1010101101;
wire [9:0] const_708_10;
assign const_708_10 = 10'b1011000100;
wire [9:0] const_990_10;
assign const_990_10 = 10'b1111011110;
wire [9:0] const_283_10;
assign const_283_10 = 10'b0100011011;
wire [9:0] const_641_10;
assign const_641_10 = 10'b1010000001;
wire [9:0] const_377_10;
assign const_377_10 = 10'b0101111001;
wire [9:0] const_160_10;
assign const_160_10 = 10'b0010100000;
wire [9:0] const_422_10;
assign const_422_10 = 10'b0110100110;
wire [9:0] const_180_10;
assign const_180_10 = 10'b0010110100;
wire [9:0] const_843_10;
assign const_843_10 = 10'b1101001011;
wire [9:0] const_704_10;
assign const_704_10 = 10'b1011000000;
wire [9:0] const_240_10;
assign const_240_10 = 10'b0011110000;
wire [9:0] const_992_10;
assign const_992_10 = 10'b1111100000;
wire [9:0] const_313_10;
assign const_313_10 = 10'b0100111001;
wire [9:0] const_545_10;
assign const_545_10 = 10'b1000100001;
wire [9:0] const_200_10;
assign const_200_10 = 10'b0011001000;
wire [9:0] const_559_10;
assign const_559_10 = 10'b1000101111;
wire [9:0] const_767_10;
assign const_767_10 = 10'b1011111111;
wire [9:0] const_551_10;
assign const_551_10 = 10'b1000100111;
wire [9:0] const_115_10;
assign const_115_10 = 10'b0001110011;
wire [9:0] const_962_10;
assign const_962_10 = 10'b1111000010;
wire [9:0] const_596_10;
assign const_596_10 = 10'b1001010100;
wire [9:0] const_98_10;
assign const_98_10 = 10'b0001100010;
wire [9:0] const_807_10;
assign const_807_10 = 10'b1100100111;
wire [9:0] const_500_10;
assign const_500_10 = 10'b0111110100;
wire [9:0] const_630_10;
assign const_630_10 = 10'b1001110110;
wire [9:0] const_451_10;
assign const_451_10 = 10'b0111000011;
wire [9:0] const_161_10;
assign const_161_10 = 10'b0010100001;
wire [9:0] const_493_10;
assign const_493_10 = 10'b0111101101;
wire [9:0] const_188_10;
assign const_188_10 = 10'b0010111100;
wire [9:0] const_544_10;
assign const_544_10 = 10'b1000100000;
wire [9:0] const_812_10;
assign const_812_10 = 10'b1100101100;
wire [9:0] const_423_10;
assign const_423_10 = 10'b0110100111;
wire [9:0] const_955_10;
assign const_955_10 = 10'b1110111011;
wire [9:0] const_906_10;
assign const_906_10 = 10'b1110001010;
wire [9:0] const_461_10;
assign const_461_10 = 10'b0111001101;
wire [9:0] const_753_10;
assign const_753_10 = 10'b1011110001;
wire [9:0] const_51_10;
assign const_51_10 = 10'b0000110011;
wire [9:0] const_856_10;
assign const_856_10 = 10'b1101011000;
wire [9:0] const_829_10;
assign const_829_10 = 10'b1100111101;
wire [9:0] const_436_10;
assign const_436_10 = 10'b0110110100;
wire [9:0] const_37_10;
assign const_37_10 = 10'b0000100101;
wire [9:0] const_408_10;
assign const_408_10 = 10'b0110011000;
wire [9:0] const_560_10;
assign const_560_10 = 10'b1000110000;
wire [9:0] const_763_10;
assign const_763_10 = 10'b1011111011;
wire [9:0] const_642_10;
assign const_642_10 = 10'b1010000010;
wire [9:0] const_419_10;
assign const_419_10 = 10'b0110100011;
wire [9:0] const_736_10;
assign const_736_10 = 10'b1011100000;
wire [9:0] const_394_10;
assign const_394_10 = 10'b0110001010;
wire [9:0] const_565_10;
assign const_565_10 = 10'b1000110101;
wire [9:0] const_538_10;
assign const_538_10 = 10'b1000011010;
wire [9:0] const_755_10;
assign const_755_10 = 10'b1011110011;
wire [9:0] const_655_10;
assign const_655_10 = 10'b1010001111;
wire [9:0] const_386_10;
assign const_386_10 = 10'b0110000010;
wire [9:0] const_201_10;
assign const_201_10 = 10'b0011001001;
wire [9:0] const_34_10;
assign const_34_10 = 10'b0000100010;
wire [9:0] const_677_10;
assign const_677_10 = 10'b1010100101;
wire [9:0] const_149_10;
assign const_149_10 = 10'b0010010101;
wire [9:0] const_588_10;
assign const_588_10 = 10'b1001001100;
wire [9:0] const_120_10;
assign const_120_10 = 10'b0001111000;
wire [9:0] const_744_10;
assign const_744_10 = 10'b1011101000;
wire [9:0] const_968_10;
assign const_968_10 = 10'b1111001000;
wire [9:0] const_626_10;
assign const_626_10 = 10'b1001110010;
wire [9:0] const_187_10;
assign const_187_10 = 10'b0010111011;
wire [9:0] const_918_10;
assign const_918_10 = 10'b1110010110;
wire [9:0] const_304_10;
assign const_304_10 = 10'b0100110000;
wire [9:0] const_5_10;
assign const_5_10 = 10'b0000000101;
wire [9:0] const_21_10;
assign const_21_10 = 10'b0000010101;
wire [9:0] const_676_10;
assign const_676_10 = 10'b1010100100;
wire [9:0] const_460_10;
assign const_460_10 = 10'b0111001100;
wire [9:0] const_153_10;
assign const_153_10 = 10'b0010011001;
wire [9:0] const_231_10;
assign const_231_10 = 10'b0011100111;
wire [9:0] const_658_10;
assign const_658_10 = 10'b1010010010;
wire [9:0] const_1014_10;
assign const_1014_10 = 10'b1111110110;
wire [9:0] const_441_10;
assign const_441_10 = 10'b0110111001;
wire [9:0] const_684_10;
assign const_684_10 = 10'b1010101100;
wire [9:0] const_443_10;
assign const_443_10 = 10'b0110111011;
wire [9:0] const_623_10;
assign const_623_10 = 10'b1001101111;
wire [9:0] const_150_10;
assign const_150_10 = 10'b0010010110;
wire [9:0] const_965_10;
assign const_965_10 = 10'b1111000101;
wire [9:0] const_432_10;
assign const_432_10 = 10'b0110110000;
wire [9:0] const_258_10;
assign const_258_10 = 10'b0100000010;
wire [9:0] const_335_10;
assign const_335_10 = 10'b0101001111;
wire [9:0] const_656_10;
assign const_656_10 = 10'b1010010000;
wire [9:0] const_546_10;
assign const_546_10 = 10'b1000100010;
wire [9:0] const_508_10;
assign const_508_10 = 10'b0111111100;
wire [9:0] const_431_10;
assign const_431_10 = 10'b0110101111;
wire [9:0] const_30_10;
assign const_30_10 = 10'b0000011110;
wire [9:0] const_840_10;
assign const_840_10 = 10'b1101001000;
wire [9:0] const_210_10;
assign const_210_10 = 10'b0011010010;
wire [9:0] const_844_10;
assign const_844_10 = 10'b1101001100;
wire [9:0] const_399_10;
assign const_399_10 = 10'b0110001111;
wire [9:0] const_391_10;
assign const_391_10 = 10'b0110000111;
wire [9:0] const_921_10;
assign const_921_10 = 10'b1110011001;
wire [9:0] const_55_10;
assign const_55_10 = 10'b0000110111;
wire [9:0] const_157_10;
assign const_157_10 = 10'b0010011101;
wire [9:0] const_657_10;
assign const_657_10 = 10'b1010010001;
wire [9:0] const_797_10;
assign const_797_10 = 10'b1100011101;
wire [9:0] const_581_10;
assign const_581_10 = 10'b1001000101;
wire [9:0] const_661_10;
assign const_661_10 = 10'b1010010101;
wire [9:0] const_699_10;
assign const_699_10 = 10'b1010111011;
wire [9:0] const_707_10;
assign const_707_10 = 10'b1011000011;
wire [9:0] const_621_10;
assign const_621_10 = 10'b1001101101;
wire [9:0] const_85_10;
assign const_85_10 = 10'b0001010101;
wire [9:0] const_574_10;
assign const_574_10 = 10'b1000111110;
wire [9:0] const_867_10;
assign const_867_10 = 10'b1101100011;
wire [9:0] const_270_10;
assign const_270_10 = 10'b0100001110;
wire [9:0] const_234_10;
assign const_234_10 = 10'b0011101010;
wire [9:0] const_311_10;
assign const_311_10 = 10'b0100110111;
wire [9:0] const_946_10;
assign const_946_10 = 10'b1110110010;
wire [9:0] const_32_10;
assign const_32_10 = 10'b0000100000;
wire [9:0] const_741_10;
assign const_741_10 = 10'b1011100101;
wire [9:0] const_524_10;
assign const_524_10 = 10'b1000001100;
wire [9:0] const_696_10;
assign const_696_10 = 10'b1010111000;
wire [9:0] const_369_10;
assign const_369_10 = 10'b0101110001;
wire [9:0] const_230_10;
assign const_230_10 = 10'b0011100110;
wire [9:0] const_532_10;
assign const_532_10 = 10'b1000010100;
wire [9:0] const_337_10;
assign const_337_10 = 10'b0101010001;
wire [9:0] const_127_10;
assign const_127_10 = 10'b0001111111;
wire [9:0] const_875_10;
assign const_875_10 = 10'b1101101011;
wire [9:0] const_207_10;
assign const_207_10 = 10'b0011001111;
wire [9:0] const_59_10;
assign const_59_10 = 10'b0000111011;

	assign comp_A1_649 = (reg_A1 <= const_649_10);
	assign comp_A2_29 = (reg_A2 <= const_29_10);
	assign comp_A3_322 = (reg_A3 <= const_322_10);
	assign comp_A4_504 = (reg_A4 <= const_504_10);
	assign comp_A5_495 = (reg_A5 <= const_495_10);
	assign comp_A6_624 = (reg_A6 <= const_624_10);
	assign comp_A7_593 = (reg_A7 <= const_593_10);
	assign comp_A1_220 = (reg_A1 <= const_220_10);
	assign comp_A4_472 = (reg_A4 <= const_472_10);
	assign comp_A8_701 = (reg_A8 <= const_701_10);
	assign comp_A9_178 = (reg_A9 <= const_178_10);
	assign comp_A91_362 = (reg_A91 <= const_362_10);
	assign comp_A92_263 = (reg_A92 <= const_263_10);
	assign comp_A93_529 = (reg_A93 <= const_529_10);
	assign comp_A94_40 = (reg_A94 <= const_40_10);
	assign comp_A7_795 = (reg_A7 <= const_795_10);
	assign comp_A95_118 = (reg_A95 <= const_118_10);
	assign comp_A3_541 = (reg_A3 <= const_541_10);
	assign comp_A8_90 = (reg_A8 <= const_90_10);
	assign comp_A96_11 = (reg_A96 <= const_11_10);
	assign comp_A97_193 = (reg_A97 <= const_193_10);
	assign comp_A98_202 = (reg_A98 <= const_202_10);
	assign comp_A99_14 = (reg_A99 <= const_14_10);
	assign comp_A2_830 = (reg_A2 <= const_830_10);
	assign comp_A991_288 = (reg_A991 <= const_288_10);
	assign comp_A992_452 = (reg_A992 <= const_452_10);
	assign comp_A95_373 = (reg_A95 <= const_373_10);
	assign comp_A8_777 = (reg_A8 <= const_777_10);
	assign comp_A93_537 = (reg_A93 <= const_537_10);
	assign comp_A99_11 = (reg_A99 <= const_11_10);
	assign comp_A95_383 = (reg_A95 <= const_383_10);
	assign comp_A993_454 = (reg_A993 <= const_454_10);
	assign comp_A992_774 = (reg_A992 <= const_774_10);
	assign comp_A994_302 = (reg_A994 <= const_302_10);
	assign comp_A995_87 = (reg_A995 <= const_87_10);
	assign comp_A98_143 = (reg_A98 <= const_143_10);
	assign comp_A996_348 = (reg_A996 <= const_348_10);
	assign comp_A997_750 = (reg_A997 <= const_750_10);
	assign comp_A1_884 = (reg_A1 <= const_884_10);
	assign comp_A997_360 = (reg_A997 <= const_360_10);
	assign comp_A998_765 = (reg_A998 <= const_765_10);
	assign comp_A8_726 = (reg_A8 <= const_726_10);
	assign comp_A999_643 = (reg_A999 <= const_643_10);
	assign comp_A3_526 = (reg_A3 <= const_526_10);
	assign comp_A7_455 = (reg_A7 <= const_455_10);
	assign comp_A9991_920 = (reg_A9991 <= const_920_10);
	assign comp_A3_300 = (reg_A3 <= const_300_10);
	assign comp_A92_262 = (reg_A92 <= const_262_10);
	assign comp_A9992_183 = (reg_A9992 <= const_183_10);
	assign comp_A991_737 = (reg_A991 <= const_737_10);
	assign comp_A97_140 = (reg_A97 <= const_140_10);
	assign comp_A9991_923 = (reg_A9991 <= const_923_10);
	assign comp_A96_873 = (reg_A96 <= const_873_10);
	assign comp_A9993_513 = (reg_A9993 <= const_513_10);
	assign comp_A4_515 = (reg_A4 <= const_515_10);
	assign comp_A9994_577 = (reg_A9994 <= const_577_10);
	assign comp_A94_46 = (reg_A94 <= const_46_10);
	assign comp_A7_341 = (reg_A7 <= const_341_10);
	assign comp_A3_687 = (reg_A3 <= const_687_10);
	assign comp_A9995_483 = (reg_A9995 <= const_483_10);
	assign comp_A9996_660 = (reg_A9996 <= const_660_10);
	assign comp_A9997_526 = (reg_A9997 <= const_526_10);
	assign comp_A9991_943 = (reg_A9991 <= const_943_10);
	assign comp_A7_561 = (reg_A7 <= const_561_10);
	assign comp_A993_276 = (reg_A993 <= const_276_10);
	assign comp_A9998_478 = (reg_A9998 <= const_478_10);
	assign comp_A92_975 = (reg_A92 <= const_975_10);
	assign comp_A1_727 = (reg_A1 <= const_727_10);
	assign comp_A7_583 = (reg_A7 <= const_583_10);
	assign comp_A995_79 = (reg_A995 <= const_79_10);
	assign comp_A97_173 = (reg_A97 <= const_173_10);
	assign comp_A993_665 = (reg_A993 <= const_665_10);
	assign comp_A9999_801 = (reg_A9999 <= const_801_10);
	assign comp_A3_536 = (reg_A3 <= const_536_10);
	assign comp_A999_620 = (reg_A999 <= const_620_10);
	assign comp_A994_700 = (reg_A994 <= const_700_10);
	assign comp_A99991_242 = (reg_A99991 <= const_242_10);
	assign comp_A994_712 = (reg_A994 <= const_712_10);
	assign comp_A99992_806 = (reg_A99992 <= const_806_10);
	assign comp_A9997_570 = (reg_A9997 <= const_570_10);
	assign comp_A99993_119 = (reg_A99993 <= const_119_10);
	assign comp_A6_670 = (reg_A6 <= const_670_10);
	assign comp_A994_338 = (reg_A994 <= const_338_10);
	assign comp_A6_635 = (reg_A6 <= const_635_10);
	assign comp_A9994_627 = (reg_A9994 <= const_627_10);
	assign comp_A1_881 = (reg_A1 <= const_881_10);
	assign comp_A4_490 = (reg_A4 <= const_490_10);
	assign comp_A92_264 = (reg_A92 <= const_264_10);
	assign comp_A2_839 = (reg_A2 <= const_839_10);
	assign comp_A991_760 = (reg_A991 <= const_760_10);
	assign comp_A993_680 = (reg_A993 <= const_680_10);
	assign comp_A99994_810 = (reg_A99994 <= const_810_10);
	assign comp_A98_974 = (reg_A98 <= const_974_10);
	assign comp_A4_350 = (reg_A4 <= const_350_10);
	assign comp_A1_738 = (reg_A1 <= const_738_10);
	assign comp_A997_319 = (reg_A997 <= const_319_10);
	assign comp_A7_411 = (reg_A7 <= const_411_10);
	assign comp_A4_400 = (reg_A4 <= const_400_10);
	assign comp_A9992_93 = (reg_A9992 <= const_93_10);
	assign comp_A99994_781 = (reg_A99994 <= const_781_10);
	assign comp_A93_726 = (reg_A93 <= const_726_10);
	assign comp_A9998_769 = (reg_A9998 <= const_769_10);
	assign comp_A7_415 = (reg_A7 <= const_415_10);
	assign comp_A9991_972 = (reg_A9991 <= const_972_10);
	assign comp_A993_608 = (reg_A993 <= const_608_10);
	assign comp_A3_284 = (reg_A3 <= const_284_10);
	assign comp_A9995_876 = (reg_A9995 <= const_876_10);
	assign comp_A9_859 = (reg_A9 <= const_859_10);
	assign comp_A9992_129 = (reg_A9992 <= const_129_10);
	assign comp_A3_102 = (reg_A3 <= const_102_10);
	assign comp_A3_79 = (reg_A3 <= const_79_10);
	assign comp_A9993_585 = (reg_A9993 <= const_585_10);
	assign comp_A3_124 = (reg_A3 <= const_124_10);
	assign comp_A91_239 = (reg_A91 <= const_239_10);
	assign comp_A93_116 = (reg_A93 <= const_116_10);
	assign comp_A9_811 = (reg_A9 <= const_811_10);
	assign comp_A3_757 = (reg_A3 <= const_757_10);
	assign comp_A99991_336 = (reg_A99991 <= const_336_10);
	assign comp_A98_66 = (reg_A98 <= const_66_10);
	assign comp_A99995_631 = (reg_A99995 <= const_631_10);
	assign comp_A999_732 = (reg_A999 <= const_732_10);
	assign comp_A9996_244 = (reg_A9996 <= const_244_10);
	assign comp_A995_167 = (reg_A995 <= const_167_10);
	assign comp_A98_171 = (reg_A98 <= const_171_10);
	assign comp_A3_981 = (reg_A3 <= const_981_10);
	assign comp_A9_827 = (reg_A9 <= const_827_10);
	assign comp_A9992_357 = (reg_A9992 <= const_357_10);
	assign comp_A4_739 = (reg_A4 <= const_739_10);
	assign comp_A2_876 = (reg_A2 <= const_876_10);
	assign comp_A99996_412 = (reg_A99996 <= const_412_10);
	assign comp_A9996_202 = (reg_A9996 <= const_202_10);
	assign comp_A9993_525 = (reg_A9993 <= const_525_10);
	assign comp_A7_666 = (reg_A7 <= const_666_10);
	assign comp_A92_519 = (reg_A92 <= const_519_10);
	assign comp_A99994_745 = (reg_A99994 <= const_745_10);
	assign comp_A998_448 = (reg_A998 <= const_448_10);
	assign comp_A9997_490 = (reg_A9997 <= const_490_10);
	assign comp_A9996_448 = (reg_A9996 <= const_448_10);
	assign comp_A997_332 = (reg_A997 <= const_332_10);
	assign comp_A4_495 = (reg_A4 <= const_495_10);
	assign comp_A94_29 = (reg_A94 <= const_29_10);
	assign comp_A7_919 = (reg_A7 <= const_919_10);
	assign comp_A99997_247 = (reg_A99997 <= const_247_10);
	assign comp_A993_764 = (reg_A993 <= const_764_10);
	assign comp_A9991_914 = (reg_A9991 <= const_914_10);
	assign comp_A96_609 = (reg_A96 <= const_609_10);
	assign comp_A9999_832 = (reg_A9999 <= const_832_10);
	assign comp_A99998_189 = (reg_A99998 <= const_189_10);
	assign comp_A996_296 = (reg_A996 <= const_296_10);
	assign comp_A99999_409 = (reg_A99999 <= const_409_10);
	assign comp_A99994_713 = (reg_A99994 <= const_713_10);
	assign comp_A993_839 = (reg_A993 <= const_839_10);
	assign comp_A99997_833 = (reg_A99997 <= const_833_10);
	assign comp_A5_327 = (reg_A5 <= const_327_10);
	assign comp_A2_894 = (reg_A2 <= const_894_10);
	assign comp_A3_587 = (reg_A3 <= const_587_10);
	assign comp_A93_629 = (reg_A93 <= const_629_10);
	assign comp_A999991_302 = (reg_A999991 <= const_302_10);
	assign comp_A99997_824 = (reg_A99997 <= const_824_10);
	assign comp_A9_155 = (reg_A9 <= const_155_10);
	assign comp_A5_170 = (reg_A5 <= const_170_10);
	assign comp_A97_991 = (reg_A97 <= const_991_10);
	assign comp_A995_114 = (reg_A995 <= const_114_10);
	assign comp_A5_586 = (reg_A5 <= const_586_10);
	assign comp_A98_162 = (reg_A98 <= const_162_10);
	assign comp_A991_728 = (reg_A991 <= const_728_10);
	assign comp_A9996_782 = (reg_A9996 <= const_782_10);
	assign comp_A99992_505 = (reg_A99992 <= const_505_10);
	assign comp_A9995_733 = (reg_A9995 <= const_733_10);
	assign comp_A9991_1016 = (reg_A9991 <= const_1016_10);
	assign comp_A9_152 = (reg_A9 <= const_152_10);
	assign comp_A5_126 = (reg_A5 <= const_126_10);
	assign comp_A999992_426 = (reg_A999992 <= const_426_10);
	assign comp_A9_784 = (reg_A9 <= const_784_10);
	assign comp_A999992_487 = (reg_A999992 <= const_487_10);
	assign comp_A92_504 = (reg_A92 <= const_504_10);
	assign comp_A9994_769 = (reg_A9994 <= const_769_10);
	assign comp_A95_435 = (reg_A95 <= const_435_10);
	assign comp_A999992_569 = (reg_A999992 <= const_569_10);
	assign comp_A1_652 = (reg_A1 <= const_652_10);
	assign comp_A991_268 = (reg_A991 <= const_268_10);
	assign comp_A99997_799 = (reg_A99997 <= const_799_10);
	assign comp_A992_599 = (reg_A992 <= const_599_10);
	assign comp_A99991_539 = (reg_A99991 <= const_539_10);
	assign comp_A98_147 = (reg_A98 <= const_147_10);
	assign comp_A7_591 = (reg_A7 <= const_591_10);
	assign comp_A997_589 = (reg_A997 <= const_589_10);
	assign comp_A97_124 = (reg_A97 <= const_124_10);
	assign comp_A996_225 = (reg_A996 <= const_225_10);
	assign comp_A97_121 = (reg_A97 <= const_121_10);
	assign comp_A99995_671 = (reg_A99995 <= const_671_10);
	assign comp_A9998_723 = (reg_A9998 <= const_723_10);
	assign comp_A999993_9 = (reg_A999993 <= const_9_10);
	assign comp_A996_92 = (reg_A996 <= const_92_10);
	assign comp_A996_222 = (reg_A996 <= const_222_10);
	assign comp_A9999_756 = (reg_A9999 <= const_756_10);
	assign comp_A95_203 = (reg_A95 <= const_203_10);
	assign comp_A997_838 = (reg_A997 <= const_838_10);
	assign comp_A5_478 = (reg_A5 <= const_478_10);
	assign comp_A99997_254 = (reg_A99997 <= const_254_10);
	assign comp_A99991_618 = (reg_A99991 <= const_618_10);
	assign comp_A91_963 = (reg_A91 <= const_963_10);
	assign comp_A9994_288 = (reg_A9994 <= const_288_10);
	assign comp_A9991_935 = (reg_A9991 <= const_935_10);
	assign comp_A99997_931 = (reg_A99997 <= const_931_10);
	assign comp_A98_151 = (reg_A98 <= const_151_10);
	assign comp_A4_486 = (reg_A4 <= const_486_10);
	assign comp_A3_232 = (reg_A3 <= const_232_10);
	assign comp_A9995_839 = (reg_A9995 <= const_839_10);
	assign comp_A7_592 = (reg_A7 <= const_592_10);
	assign comp_A3_286 = (reg_A3 <= const_286_10);
	assign comp_A99999_486 = (reg_A99999 <= const_486_10);
	assign comp_A9991_932 = (reg_A9991 <= const_932_10);
	assign comp_A996_372 = (reg_A996 <= const_372_10);
	assign comp_A9_156 = (reg_A9 <= const_156_10);
	assign comp_A7_804 = (reg_A7 <= const_804_10);
	assign comp_A6_255 = (reg_A6 <= const_255_10);
	assign comp_A99991_344 = (reg_A99991 <= const_344_10);
	assign comp_A8_757 = (reg_A8 <= const_757_10);
	assign comp_A993_555 = (reg_A993 <= const_555_10);
	assign comp_A999994_442 = (reg_A999994 <= const_442_10);
	assign comp_A99992_671 = (reg_A99992 <= const_671_10);
	assign comp_A991_479 = (reg_A991 <= const_479_10);
	assign comp_A97_610 = (reg_A97 <= const_610_10);
	assign comp_A999991_570 = (reg_A999991 <= const_570_10);
	assign comp_A9_816 = (reg_A9 <= const_816_10);
	assign comp_A3_80 = (reg_A3 <= const_80_10);
	assign comp_A8_822 = (reg_A8 <= const_822_10);
	assign comp_A998_424 = (reg_A998 <= const_424_10);
	assign comp_A999993_8 = (reg_A999993 <= const_8_10);
	assign comp_A9992_421 = (reg_A9992 <= const_421_10);
	assign comp_A99999_549 = (reg_A99999 <= const_549_10);
	assign comp_A9993_307 = (reg_A9993 <= const_307_10);
	assign comp_A9996_562 = (reg_A9996 <= const_562_10);
	assign comp_A996_271 = (reg_A996 <= const_271_10);
	assign comp_A992_400 = (reg_A992 <= const_400_10);
	assign comp_A94_31 = (reg_A94 <= const_31_10);
	assign comp_A99_8 = (reg_A99 <= const_8_10);
	assign comp_A3_54 = (reg_A3 <= const_54_10);
	assign comp_A2_872 = (reg_A2 <= const_872_10);
	assign comp_A92_972 = (reg_A92 <= const_972_10);
	assign comp_A3_272 = (reg_A3 <= const_272_10);
	assign comp_A999995_1015 = (reg_A999995 <= const_1015_10);
	assign comp_A7_605 = (reg_A7 <= const_605_10);
	assign comp_A9993_295 = (reg_A9993 <= const_295_10);
	assign comp_A991_531 = (reg_A991 <= const_531_10);
	assign comp_A993_317 = (reg_A993 <= const_317_10);
	assign comp_A991_869 = (reg_A991 <= const_869_10);
	assign comp_A94_50 = (reg_A94 <= const_50_10);
	assign comp_A99994_178 = (reg_A99994 <= const_178_10);
	assign comp_A8_786 = (reg_A8 <= const_786_10);
	assign comp_A3_407 = (reg_A3 <= const_407_10);
	assign comp_A6_722 = (reg_A6 <= const_722_10);
	assign comp_A99999_735 = (reg_A99999 <= const_735_10);
	assign comp_A92_259 = (reg_A92 <= const_259_10);
	assign comp_A999996_390 = (reg_A999996 <= const_390_10);
	assign comp_A2_901 = (reg_A2 <= const_901_10);
	assign comp_A992_675 = (reg_A992 <= const_675_10);
	assign comp_A9_821 = (reg_A9 <= const_821_10);
	assign comp_A92_503 = (reg_A92 <= const_503_10);
	assign comp_A8_536 = (reg_A8 <= const_536_10);
	assign comp_A2_124 = (reg_A2 <= const_124_10);
	assign comp_A92_250 = (reg_A92 <= const_250_10);
	assign comp_A95_497 = (reg_A95 <= const_497_10);
	assign comp_A6_406 = (reg_A6 <= const_406_10);
	assign comp_A9991_948 = (reg_A9991 <= const_948_10);
	assign comp_A9999_819 = (reg_A9999 <= const_819_10);
	assign comp_A3_535 = (reg_A3 <= const_535_10);
	assign comp_A998_805 = (reg_A998 <= const_805_10);
	assign comp_A92_995 = (reg_A92 <= const_995_10);
	assign comp_A9996_600 = (reg_A9996 <= const_600_10);
	assign comp_A6_606 = (reg_A6 <= const_606_10);
	assign comp_A996_353 = (reg_A996 <= const_353_10);
	assign comp_A99994_600 = (reg_A99994 <= const_600_10);
	assign comp_A99991_286 = (reg_A99991 <= const_286_10);
	assign comp_A996_340 = (reg_A996 <= const_340_10);
	assign comp_A998_414 = (reg_A998 <= const_414_10);
	assign comp_A996_331 = (reg_A996 <= const_331_10);
	assign comp_A994_640 = (reg_A994 <= const_640_10);
	assign comp_A999_714 = (reg_A999 <= const_714_10);
	assign comp_A3_233 = (reg_A3 <= const_233_10);
	assign comp_A9_805 = (reg_A9 <= const_805_10);
	assign comp_A8_540 = (reg_A8 <= const_540_10);
	assign comp_A99996_575 = (reg_A99996 <= const_575_10);
	assign comp_A993_982 = (reg_A993 <= const_982_10);
	assign comp_A9993_530 = (reg_A9993 <= const_530_10);
	assign comp_A994_475 = (reg_A994 <= const_475_10);
	assign comp_A996_332 = (reg_A996 <= const_332_10);
	assign comp_A4_484 = (reg_A4 <= const_484_10);
	assign comp_A98_325 = (reg_A98 <= const_325_10);
	assign comp_A993_659 = (reg_A993 <= const_659_10);
	assign comp_A2_602 = (reg_A2 <= const_602_10);
	assign comp_A92_505 = (reg_A92 <= const_505_10);
	assign comp_A99999_58 = (reg_A99999 <= const_58_10);
	assign comp_A9992_123 = (reg_A9992 <= const_123_10);
	assign comp_A999992_527 = (reg_A999992 <= const_527_10);
	assign comp_A9996_758 = (reg_A9996 <= const_758_10);
	assign comp_A997_428 = (reg_A997 <= const_428_10);
	assign comp_A3_515 = (reg_A3 <= const_515_10);
	assign comp_A992_389 = (reg_A992 <= const_389_10);
	assign comp_A93_513 = (reg_A93 <= const_513_10);
	assign comp_A99999_558 = (reg_A99999 <= const_558_10);
	assign comp_A9992_429 = (reg_A9992 <= const_429_10);
	assign comp_A993_440 = (reg_A993 <= const_440_10);
	assign comp_A99996_766 = (reg_A99996 <= const_766_10);
	assign comp_A999991_485 = (reg_A999991 <= const_485_10);
	assign comp_A9991_1009 = (reg_A9991 <= const_1009_10);
	assign comp_A99999_594 = (reg_A99999 <= const_594_10);
	assign comp_A993_492 = (reg_A993 <= const_492_10);
	assign comp_A96_754 = (reg_A96 <= const_754_10);
	assign comp_A993_321 = (reg_A993 <= const_321_10);
	assign comp_A999_712 = (reg_A999 <= const_712_10);
	assign comp_A997_421 = (reg_A997 <= const_421_10);
	assign comp_A9999_805 = (reg_A9999 <= const_805_10);
	assign comp_A995_343 = (reg_A995 <= const_343_10);
	assign comp_A9996_570 = (reg_A9996 <= const_570_10);
	assign comp_A5_653 = (reg_A5 <= const_653_10);
	assign comp_A4_445 = (reg_A4 <= const_445_10);
	assign comp_A99995_511 = (reg_A99995 <= const_511_10);
	assign comp_A99991_185 = (reg_A99991 <= const_185_10);
	assign comp_A99999_517 = (reg_A99999 <= const_517_10);
	assign comp_A8_334 = (reg_A8 <= const_334_10);
	assign comp_A9996_737 = (reg_A9996 <= const_737_10);
	assign comp_A9_845 = (reg_A9 <= const_845_10);
	assign comp_A997_339 = (reg_A997 <= const_339_10);
	assign comp_A997_243 = (reg_A997 <= const_243_10);
	assign comp_A993_683 = (reg_A993 <= const_683_10);
	assign comp_A994_543 = (reg_A994 <= const_543_10);
	assign comp_A99_13 = (reg_A99 <= const_13_10);
	assign comp_A2_22 = (reg_A2 <= const_22_10);
	assign comp_A96_818 = (reg_A96 <= const_818_10);
	assign comp_A3_350 = (reg_A3 <= const_350_10);
	assign comp_A992_528 = (reg_A992 <= const_528_10);
	assign comp_A96_271 = (reg_A96 <= const_271_10);
	assign comp_A994_365 = (reg_A994 <= const_365_10);
	assign comp_A999991_372 = (reg_A999991 <= const_372_10);
	assign comp_A99999_168 = (reg_A99999 <= const_168_10);
	assign comp_A95_430 = (reg_A95 <= const_430_10);
	assign comp_A8_398 = (reg_A8 <= const_398_10);
	assign comp_A994_484 = (reg_A994 <= const_484_10);
	assign comp_A999997_1009 = (reg_A999997 <= const_1009_10);
	assign comp_A3_415 = (reg_A3 <= const_415_10);
	assign comp_A97_174 = (reg_A97 <= const_174_10);
	assign comp_A997_549 = (reg_A997 <= const_549_10);
	assign comp_A999996_427 = (reg_A999996 <= const_427_10);
	assign comp_A3_381 = (reg_A3 <= const_381_10);
	assign comp_A997_496 = (reg_A997 <= const_496_10);
	assign comp_A995_61 = (reg_A995 <= const_61_10);
	assign comp_A99_15 = (reg_A99 <= const_15_10);
	assign comp_A99_18 = (reg_A99 <= const_18_10);
	assign comp_A992_721 = (reg_A992 <= const_721_10);
	assign comp_A6_474 = (reg_A6 <= const_474_10);
	assign comp_A95_345 = (reg_A95 <= const_345_10);
	assign comp_A2_860 = (reg_A2 <= const_860_10);
	assign comp_A9_853 = (reg_A9 <= const_853_10);
	assign comp_A93_136 = (reg_A93 <= const_136_10);
	assign comp_A991_746 = (reg_A991 <= const_746_10);
	assign comp_A2_320 = (reg_A2 <= const_320_10);
	assign comp_A97_182 = (reg_A97 <= const_182_10);
	assign comp_A91_383 = (reg_A91 <= const_383_10);
	assign comp_A6_485 = (reg_A6 <= const_485_10);
	assign comp_A99995_471 = (reg_A99995 <= const_471_10);
	assign comp_A93_516 = (reg_A93 <= const_516_10);
	assign comp_A99992_501 = (reg_A99992 <= const_501_10);
	assign comp_A2_920 = (reg_A2 <= const_920_10);
	assign comp_A9991_961 = (reg_A9991 <= const_961_10);
	assign comp_A999996_360 = (reg_A999996 <= const_360_10);
	assign comp_A996_350 = (reg_A996 <= const_350_10);
	assign comp_A991_868 = (reg_A991 <= const_868_10);
	assign comp_A992_266 = (reg_A992 <= const_266_10);
	assign comp_A95_312 = (reg_A95 <= const_312_10);
	assign comp_A96_171 = (reg_A96 <= const_171_10);
	assign comp_A98_61 = (reg_A98 <= const_61_10);
	assign comp_A9994_693 = (reg_A9994 <= const_693_10);
	assign comp_A994_378 = (reg_A994 <= const_378_10);
	assign comp_A99991_182 = (reg_A99991 <= const_182_10);
	assign comp_A8_718 = (reg_A8 <= const_718_10);
	assign comp_A3_428 = (reg_A3 <= const_428_10);
	assign comp_A99996_862 = (reg_A99996 <= const_862_10);
	assign comp_A9993_327 = (reg_A9993 <= const_327_10);
	assign comp_A995_537 = (reg_A995 <= const_537_10);
	assign comp_A9_832 = (reg_A9 <= const_832_10);
	assign comp_A6_442 = (reg_A6 <= const_442_10);
	assign comp_A999996_428 = (reg_A999996 <= const_428_10);
	assign comp_A94_58 = (reg_A94 <= const_58_10);
	assign comp_A997_521 = (reg_A997 <= const_521_10);
	assign comp_A996_360 = (reg_A996 <= const_360_10);
	assign comp_A99992_503 = (reg_A99992 <= const_503_10);
	assign comp_A999994_457 = (reg_A999994 <= const_457_10);
	assign comp_A99992_710 = (reg_A99992 <= const_710_10);
	assign comp_A99991_366 = (reg_A99991 <= const_366_10);
	assign comp_A993_286 = (reg_A993 <= const_286_10);
	assign comp_A999_567 = (reg_A999 <= const_567_10);
	assign comp_A99996_858 = (reg_A99996 <= const_858_10);
	assign comp_A5_316 = (reg_A5 <= const_316_10);
	assign comp_A995_299 = (reg_A995 <= const_299_10);
	assign comp_A991_852 = (reg_A991 <= const_852_10);
	assign comp_A94_49 = (reg_A94 <= const_49_10);
	assign comp_A9992_105 = (reg_A9992 <= const_105_10);
	assign comp_A92_247 = (reg_A92 <= const_247_10);
	assign comp_A98_68 = (reg_A98 <= const_68_10);
	assign comp_A99995_519 = (reg_A99995 <= const_519_10);
	assign comp_A92_989 = (reg_A92 <= const_989_10);
	assign comp_A3_285 = (reg_A3 <= const_285_10);
	assign comp_A94_42 = (reg_A94 <= const_42_10);
	assign comp_A97_400 = (reg_A97 <= const_400_10);
	assign comp_A3_209 = (reg_A3 <= const_209_10);
	assign comp_A8_381 = (reg_A8 <= const_381_10);
	assign comp_A99_19 = (reg_A99 <= const_19_10);
	assign comp_A999997_1011 = (reg_A999997 <= const_1011_10);
	assign comp_A92_815 = (reg_A92 <= const_815_10);
	assign comp_A94_33 = (reg_A94 <= const_33_10);
	assign comp_A9991_937 = (reg_A9991 <= const_937_10);
	assign comp_A998_499 = (reg_A998 <= const_499_10);
	assign comp_A1_554 = (reg_A1 <= const_554_10);
	assign comp_A999994_662 = (reg_A999994 <= const_662_10);
	assign comp_A5_562 = (reg_A5 <= const_562_10);
	assign comp_A9997_669 = (reg_A9997 <= const_669_10);
	assign comp_A997_477 = (reg_A997 <= const_477_10);
	assign comp_A9991_973 = (reg_A9991 <= const_973_10);
	assign comp_A9999_248 = (reg_A9999 <= const_248_10);
	assign comp_A996_245 = (reg_A996 <= const_245_10);
	assign comp_A98_1019 = (reg_A98 <= const_1019_10);
	assign comp_A3_112 = (reg_A3 <= const_112_10);
	assign comp_A994_355 = (reg_A994 <= const_355_10);
	assign comp_A993_548 = (reg_A993 <= const_548_10);
	assign comp_A9991_817 = (reg_A9991 <= const_817_10);
	assign comp_A92_246 = (reg_A92 <= const_246_10);
	assign comp_A3_27 = (reg_A3 <= const_27_10);
	assign comp_A8_810 = (reg_A8 <= const_810_10);
	assign comp_A99994_682 = (reg_A99994 <= const_682_10);
	assign comp_A993_612 = (reg_A993 <= const_612_10);
	assign comp_A9992_99 = (reg_A9992 <= const_99_10);
	assign comp_A9996_610 = (reg_A9996 <= const_610_10);
	assign comp_A997_620 = (reg_A997 <= const_620_10);
	assign comp_A994_477 = (reg_A994 <= const_477_10);
	assign comp_A9999_293 = (reg_A9999 <= const_293_10);
	assign comp_A8_404 = (reg_A8 <= const_404_10);
	assign comp_A996_318 = (reg_A996 <= const_318_10);
	assign comp_A95_274 = (reg_A95 <= const_274_10);
	assign comp_A1_601 = (reg_A1 <= const_601_10);
	assign comp_A92_562 = (reg_A92 <= const_562_10);
	assign comp_A99997_252 = (reg_A99997 <= const_252_10);
	assign comp_A9996_694 = (reg_A9996 <= const_694_10);
	assign comp_A3_305 = (reg_A3 <= const_305_10);
	assign comp_A997_334 = (reg_A997 <= const_334_10);
	assign comp_A999994_507 = (reg_A999994 <= const_507_10);
	assign comp_A99993_647 = (reg_A99993 <= const_647_10);
	assign comp_A992_308 = (reg_A992 <= const_308_10);
	assign comp_A99992_810 = (reg_A99992 <= const_810_10);
	assign comp_A9993_652 = (reg_A9993 <= const_652_10);
	assign comp_A997_403 = (reg_A997 <= const_403_10);
	assign comp_A93_651 = (reg_A93 <= const_651_10);
	assign comp_A999991_306 = (reg_A999991 <= const_306_10);
	assign comp_A991_720 = (reg_A991 <= const_720_10);
	assign comp_A9992_107 = (reg_A9992 <= const_107_10);
	assign comp_A9_851 = (reg_A9 <= const_851_10);
	assign comp_A9992_103 = (reg_A9992 <= const_103_10);
	assign comp_A2_869 = (reg_A2 <= const_869_10);
	assign comp_A997_578 = (reg_A997 <= const_578_10);
	assign comp_A998_302 = (reg_A998 <= const_302_10);
	assign comp_A99991_660 = (reg_A99991 <= const_660_10);
	assign comp_A6_644 = (reg_A6 <= const_644_10);
	assign comp_A2_285 = (reg_A2 <= const_285_10);
	assign comp_A995_202 = (reg_A995 <= const_202_10);
	assign comp_A8_818 = (reg_A8 <= const_818_10);
	assign comp_A999995_1012 = (reg_A999995 <= const_1012_10);
	assign comp_A997_956 = (reg_A997 <= const_956_10);
	assign comp_A999992_388 = (reg_A999992 <= const_388_10);
	assign comp_A93_687 = (reg_A93 <= const_687_10);
	assign comp_A999995_1008 = (reg_A999995 <= const_1008_10);
	assign comp_A996_292 = (reg_A996 <= const_292_10);
	assign comp_A991_250 = (reg_A991 <= const_250_10);
	assign comp_A95_354 = (reg_A95 <= const_354_10);
	assign comp_A9994_711 = (reg_A9994 <= const_711_10);
	assign comp_A9994_295 = (reg_A9994 <= const_295_10);
	assign comp_A5_505 = (reg_A5 <= const_505_10);
	assign comp_A94_35 = (reg_A94 <= const_35_10);
	assign comp_A999994_547 = (reg_A999994 <= const_547_10);
	assign comp_A9993_685 = (reg_A9993 <= const_685_10);
	assign comp_A93_718 = (reg_A93 <= const_718_10);
	assign comp_A9991_956 = (reg_A9991 <= const_956_10);
	assign comp_A993_484 = (reg_A993 <= const_484_10);
	assign comp_A1_708 = (reg_A1 <= const_708_10);
	assign comp_A9991_990 = (reg_A9991 <= const_990_10);
	assign comp_A3_283 = (reg_A3 <= const_283_10);
	assign comp_A998_641 = (reg_A998 <= const_641_10);
	assign comp_A92_377 = (reg_A92 <= const_377_10);
	assign comp_A99994_383 = (reg_A99994 <= const_383_10);
	assign comp_A999992_484 = (reg_A999992 <= const_484_10);
	assign comp_A9_160 = (reg_A9 <= const_160_10);
	assign comp_A997_422 = (reg_A997 <= const_422_10);
	assign comp_A2_862 = (reg_A2 <= const_862_10);
	assign comp_A96_180 = (reg_A96 <= const_180_10);
	assign comp_A99997_843 = (reg_A99997 <= const_843_10);
	assign comp_A9994_704 = (reg_A9994 <= const_704_10);
	assign comp_A98_240 = (reg_A98 <= const_240_10);
	assign comp_A3_992 = (reg_A3 <= const_992_10);
	assign comp_A9994_881 = (reg_A9994 <= const_881_10);
	assign comp_A2_827 = (reg_A2 <= const_827_10);
	assign comp_A999997_1012 = (reg_A999997 <= const_1012_10);
	assign comp_A994_549 = (reg_A994 <= const_549_10);
	assign comp_A97_171 = (reg_A97 <= const_171_10);
	assign comp_A9993_313 = (reg_A9993 <= const_313_10);
	assign comp_A4_545 = (reg_A4 <= const_545_10);
	assign comp_A996_200 = (reg_A996 <= const_200_10);
	assign comp_A3_247 = (reg_A3 <= const_247_10);
	assign comp_A995_185 = (reg_A995 <= const_185_10);
	assign comp_A998_559 = (reg_A998 <= const_559_10);
	assign comp_A9999_767 = (reg_A9999 <= const_767_10);
	assign comp_A99996_551 = (reg_A99996 <= const_551_10);
	assign comp_A6_701 = (reg_A6 <= const_701_10);
	assign comp_A992_817 = (reg_A992 <= const_817_10);
	assign comp_A93_115 = (reg_A93 <= const_115_10);
	assign comp_A9991_962 = (reg_A9991 <= const_962_10);
	assign comp_A99993_596 = (reg_A99993 <= const_596_10);
	assign comp_A93_98 = (reg_A93 <= const_98_10);
	assign comp_A99994_807 = (reg_A99994 <= const_807_10);
	assign comp_A96_264 = (reg_A96 <= const_264_10);
	assign comp_A92_500 = (reg_A92 <= const_500_10);
	assign comp_A9996_693 = (reg_A9996 <= const_693_10);
	assign comp_A99993_630 = (reg_A99993 <= const_630_10);
	assign comp_A99996_513 = (reg_A99996 <= const_513_10);
	assign comp_A997_451 = (reg_A997 <= const_451_10);
	assign comp_A9992_161 = (reg_A9992 <= const_161_10);
	assign comp_A2_114 = (reg_A2 <= const_114_10);
	assign comp_A995_493 = (reg_A995 <= const_493_10);
	assign comp_A99996_188 = (reg_A99996 <= const_188_10);
	assign comp_A3_116 = (reg_A3 <= const_116_10);
	assign comp_A99996_839 = (reg_A99996 <= const_839_10);
	assign comp_A2_9 = (reg_A2 <= const_9_10);
	assign comp_A93_544 = (reg_A93 <= const_544_10);
	assign comp_A3_812 = (reg_A3 <= const_812_10);
	assign comp_A997_373 = (reg_A997 <= const_373_10);
	assign comp_A99999_423 = (reg_A99999 <= const_423_10);
	assign comp_A9991_955 = (reg_A9991 <= const_955_10);
	assign comp_A9998_906 = (reg_A9998 <= const_906_10);
	assign comp_A999996_461 = (reg_A999996 <= const_461_10);
	assign comp_A999_585 = (reg_A999 <= const_585_10);
	assign comp_A5_753 = (reg_A5 <= const_753_10);
	assign comp_A99993_51 = (reg_A99993 <= const_51_10);
	assign comp_A92_255 = (reg_A92 <= const_255_10);
	assign comp_A7_856 = (reg_A7 <= const_856_10);
	assign comp_A9_829 = (reg_A9 <= const_829_10);
	assign comp_A99995_559 = (reg_A99995 <= const_559_10);
	assign comp_A2_33 = (reg_A2 <= const_33_10);
	assign comp_A99999_545 = (reg_A99999 <= const_545_10);
	assign comp_A9992_436 = (reg_A9992 <= const_436_10);
	assign comp_A997_666 = (reg_A997 <= const_666_10);
	assign comp_A94_37 = (reg_A94 <= const_37_10);
	assign comp_A9991_1011 = (reg_A9991 <= const_1011_10);
	assign comp_A99991_408 = (reg_A99991 <= const_408_10);
	assign comp_A996_343 = (reg_A996 <= const_343_10);
	assign comp_A9999_560 = (reg_A9999 <= const_560_10);
	assign comp_A996_263 = (reg_A996 <= const_263_10);
	assign comp_A9996_763 = (reg_A9996 <= const_763_10);
	assign comp_A99992_660 = (reg_A99992 <= const_660_10);
	assign comp_A1_642 = (reg_A1 <= const_642_10);
	assign comp_A9999_419 = (reg_A9999 <= const_419_10);
	assign comp_A7_643 = (reg_A7 <= const_643_10);
	assign comp_A99992_736 = (reg_A99992 <= const_736_10);
	assign comp_A9_61 = (reg_A9 <= const_61_10);
	assign comp_A6_394 = (reg_A6 <= const_394_10);
	assign comp_A99999_406 = (reg_A99999 <= const_406_10);
	assign comp_A3_565 = (reg_A3 <= const_565_10);
	assign comp_A997_381 = (reg_A997 <= const_381_10);
	assign comp_A99992_538 = (reg_A99992 <= const_538_10);
	assign comp_A99994_755 = (reg_A99994 <= const_755_10);
	assign comp_A8_484 = (reg_A8 <= const_484_10);
	assign comp_A99992_655 = (reg_A99992 <= const_655_10);
	assign comp_A991_451 = (reg_A991 <= const_451_10);
	assign comp_A99995_531 = (reg_A99995 <= const_531_10);
	assign comp_A3_386 = (reg_A3 <= const_386_10);
	assign comp_A9998_389 = (reg_A9998 <= const_389_10);
	assign comp_A994_390 = (reg_A994 <= const_390_10);
	assign comp_A97_201 = (reg_A97 <= const_201_10);
	assign comp_A3_750 = (reg_A3 <= const_750_10);
	assign comp_A995_34 = (reg_A995 <= const_34_10);
	assign comp_A994_677 = (reg_A994 <= const_677_10);
	assign comp_A93_720 = (reg_A93 <= const_720_10);
	assign comp_A99997_149 = (reg_A99997 <= const_149_10);
	assign comp_A3_588 = (reg_A3 <= const_588_10);
	assign comp_A98_120 = (reg_A98 <= const_120_10);
	assign comp_A9_151 = (reg_A9 <= const_151_10);
	assign comp_A996_244 = (reg_A996 <= const_244_10);
	assign comp_A9999_786 = (reg_A9999 <= const_786_10);
	assign comp_A99992_744 = (reg_A99992 <= const_744_10);
	assign comp_A97_968 = (reg_A97 <= const_968_10);
	assign comp_A9993_626 = (reg_A9993 <= const_626_10);
	assign comp_A99998_187 = (reg_A99998 <= const_187_10);
	assign comp_A99994_612 = (reg_A99994 <= const_612_10);
	assign comp_A9991_982 = (reg_A9991 <= const_982_10);
	assign comp_A2_918 = (reg_A2 <= const_918_10);
	assign comp_A996_304 = (reg_A996 <= const_304_10);
	assign comp_A99_5 = (reg_A99 <= const_5_10);
	assign comp_A9991_693 = (reg_A9991 <= const_693_10);
	assign comp_A99_21 = (reg_A99 <= const_21_10);
	assign comp_A9991_931 = (reg_A9991 <= const_931_10);
	assign comp_A3_103 = (reg_A3 <= const_103_10);
	assign comp_A998_676 = (reg_A998 <= const_676_10);
	assign comp_A9_486 = (reg_A9 <= const_486_10);
	assign comp_A92_528 = (reg_A92 <= const_528_10);
	assign comp_A7_460 = (reg_A7 <= const_460_10);
	assign comp_A999994_411 = (reg_A999994 <= const_411_10);
	assign comp_A93_722 = (reg_A93 <= const_722_10);
	assign comp_A98_153 = (reg_A98 <= const_153_10);
	assign comp_A996_231 = (reg_A996 <= const_231_10);
	assign comp_A999_516 = (reg_A999 <= const_516_10);
	assign comp_A991_373 = (reg_A991 <= const_373_10);
	assign comp_A9993_658 = (reg_A9993 <= const_658_10);
	assign comp_A999992_474 = (reg_A999992 <= const_474_10);
	assign comp_A999995_1014 = (reg_A999995 <= const_1014_10);
	assign comp_A9995_441 = (reg_A9995 <= const_441_10);
	assign comp_A996_327 = (reg_A996 <= const_327_10);
	assign comp_A1_684 = (reg_A1 <= const_684_10);
	assign comp_A99999_443 = (reg_A99999 <= const_443_10);
	assign comp_A9996_623 = (reg_A9996 <= const_623_10);
	assign comp_A9_150 = (reg_A9 <= const_150_10);
	assign comp_A997_713 = (reg_A997 <= const_713_10);
	assign comp_A9991_965 = (reg_A9991 <= const_965_10);
	assign comp_A999992_432 = (reg_A999992 <= const_432_10);
	assign comp_A999996_726 = (reg_A999996 <= const_726_10);
	assign comp_A993_258 = (reg_A993 <= const_258_10);
	assign comp_A8_335 = (reg_A8 <= const_335_10);
	assign comp_A999_656 = (reg_A999 <= const_656_10);
	assign comp_A991_735 = (reg_A991 <= const_735_10);
	assign comp_A996_203 = (reg_A996 <= const_203_10);
	assign comp_A93_546 = (reg_A93 <= const_546_10);
	assign comp_A99996_508 = (reg_A99996 <= const_508_10);
	assign comp_A99996_263 = (reg_A99996 <= const_263_10);
	assign comp_A9996_431 = (reg_A9996 <= const_431_10);
	assign comp_A96_22 = (reg_A96 <= const_22_10);
	assign comp_A94_30 = (reg_A94 <= const_30_10);
	assign comp_A999_711 = (reg_A999 <= const_711_10);
	assign comp_A9_840 = (reg_A9 <= const_840_10);
	assign comp_A91_210 = (reg_A91 <= const_210_10);
	assign comp_A9997_587 = (reg_A9997 <= const_587_10);
	assign comp_A2_713 = (reg_A2 <= const_713_10);
	assign comp_A999996_685 = (reg_A999996 <= const_685_10);
	assign comp_A2_844 = (reg_A2 <= const_844_10);
	assign comp_A997_399 = (reg_A997 <= const_399_10);
	assign comp_A9993_561 = (reg_A9993 <= const_561_10);
	assign comp_A991_391 = (reg_A991 <= const_391_10);
	assign comp_A6_286 = (reg_A6 <= const_286_10);
	assign comp_A99992_711 = (reg_A99992 <= const_711_10);
	assign comp_A9991_921 = (reg_A9991 <= const_921_10);
	assign comp_A3_55 = (reg_A3 <= const_55_10);
	assign comp_A9_157 = (reg_A9 <= const_157_10);
	assign comp_A8_657 = (reg_A8 <= const_657_10);
	assign comp_A99994_586 = (reg_A99994 <= const_586_10);
	assign comp_A991_797 = (reg_A991 <= const_797_10);
	assign comp_A997_394 = (reg_A997 <= const_394_10);
	assign comp_A96_766 = (reg_A96 <= const_766_10);
	assign comp_A9993_581 = (reg_A9993 <= const_581_10);
	assign comp_A9998_661 = (reg_A9998 <= const_661_10);
	assign comp_A99993_699 = (reg_A99993 <= const_699_10);
	assign comp_A9996_707 = (reg_A9996 <= const_707_10);
	assign comp_A99997_955 = (reg_A99997 <= const_955_10);
	assign comp_A991_647 = (reg_A991 <= const_647_10);
	assign comp_A996_185 = (reg_A996 <= const_185_10);
	assign comp_A999992_536 = (reg_A999992 <= const_536_10);
	assign comp_A93_92 = (reg_A93 <= const_92_10);
	assign comp_A1_581 = (reg_A1 <= const_581_10);
	assign comp_A991_486 = (reg_A991 <= const_486_10);
	assign comp_A993_621 = (reg_A993 <= const_621_10);
	assign comp_A999992_339 = (reg_A999992 <= const_339_10);
	assign comp_A7_767 = (reg_A7 <= const_767_10);
	assign comp_A99993_85 = (reg_A99993 <= const_85_10);
	assign comp_A92_574 = (reg_A92 <= const_574_10);
	assign comp_A3_867 = (reg_A3 <= const_867_10);
	assign comp_A98_270 = (reg_A98 <= const_270_10);
	assign comp_A93_119 = (reg_A93 <= const_119_10);
	assign comp_A992_234 = (reg_A992 <= const_234_10);
	assign comp_A92_992 = (reg_A92 <= const_992_10);
	assign comp_A991_644 = (reg_A991 <= const_644_10);
	assign comp_A3_662 = (reg_A3 <= const_662_10);
	assign comp_A996_311 = (reg_A996 <= const_311_10);
	assign comp_A994_457 = (reg_A994 <= const_457_10);
	assign comp_A9993_539 = (reg_A9993 <= const_539_10);
	assign comp_A99997_946 = (reg_A99997 <= const_946_10);
	assign comp_A997_299 = (reg_A997 <= const_299_10);
	assign comp_A99992_670 = (reg_A99992 <= const_670_10);
	assign comp_A94_32 = (reg_A94 <= const_32_10);
	assign comp_A1_741 = (reg_A1 <= const_741_10);
	assign comp_A994_524 = (reg_A994 <= const_524_10);
	assign comp_A9997_340 = (reg_A9997 <= const_340_10);
	assign comp_A997_696 = (reg_A997 <= const_696_10);
	assign comp_A99994_727 = (reg_A99994 <= const_727_10);
	assign comp_A994_644 = (reg_A994 <= const_644_10);
	assign comp_A996_369 = (reg_A996 <= const_369_10);
	assign comp_A9991_995 = (reg_A9991 <= const_995_10);
	assign comp_A5_492 = (reg_A5 <= const_492_10);
	assign comp_A998_230 = (reg_A998 <= const_230_10);
	assign comp_A93_532 = (reg_A93 <= const_532_10);
	assign comp_A999_337 = (reg_A999 <= const_337_10);
	assign comp_A95_388 = (reg_A95 <= const_388_10);
	assign comp_A3_127 = (reg_A3 <= const_127_10);
	assign comp_A6_452 = (reg_A6 <= const_452_10);
	assign comp_A4_332 = (reg_A4 <= const_332_10);
	assign comp_A999996_581 = (reg_A999996 <= const_581_10);
	assign comp_A8_875 = (reg_A8 <= const_875_10);
	assign comp_A97_207 = (reg_A97 <= const_207_10);
	assign comp_A9993_671 = (reg_A9993 <= const_671_10);
	assign comp_A9999_59 = (reg_A9999 <= const_59_10);
	assign comp_A991_777 = (reg_A991 <= const_777_10);
	assign comp_A9991_699 = (reg_A9991 <= const_699_10);
endmodule


module ANDS(
comp_A1_649, comp_A2_29, comp_A3_322, comp_A4_504, comp_A5_495, comp_A6_624, comp_A7_593, comp_A1_220, comp_A4_472, comp_A8_701, comp_A9_178, comp_A91_362, comp_A92_263, comp_A93_529, comp_A94_40, comp_A7_795, comp_A95_118, comp_A3_541, comp_A8_90, comp_A96_11, comp_A97_193, comp_A98_202, comp_A99_14, comp_A2_830, comp_A991_288, comp_A992_452, comp_A95_373, comp_A8_777, comp_A93_537, comp_A99_11, comp_A95_383, comp_A993_454, comp_A992_774, comp_A994_302, comp_A995_87, comp_A98_143, comp_A996_348, comp_A997_750, comp_A1_884, comp_A997_360, comp_A998_765, comp_A8_726, comp_A999_643, comp_A3_526, comp_A7_455, comp_A9991_920, comp_A3_300, comp_A92_262, comp_A9992_183, comp_A991_737, comp_A97_140, comp_A9991_923, comp_A96_873, comp_A9993_513, comp_A4_515, comp_A9994_577, comp_A94_46, comp_A7_341, comp_A3_687, comp_A9995_483, comp_A9996_660, comp_A9997_526, comp_A9991_943, comp_A7_561, comp_A993_276, comp_A9998_478, comp_A92_975, comp_A1_727, comp_A7_583, comp_A995_79, comp_A97_173, comp_A993_665, comp_A9999_801, comp_A3_536, comp_A999_620, comp_A994_700, comp_A99991_242, comp_A994_712, comp_A99992_806, comp_A9997_570, comp_A99993_119, comp_A6_670, comp_A994_338, comp_A6_635, comp_A9994_627, comp_A1_881, comp_A4_490, comp_A92_264, comp_A2_839, comp_A991_760, comp_A993_680, comp_A99994_810, comp_A98_974, comp_A4_350, comp_A1_738, comp_A997_319, comp_A7_411, comp_A4_400, comp_A9992_93, comp_A99994_781, comp_A93_726, comp_A9998_769, comp_A7_415, comp_A9991_972, comp_A993_608, comp_A3_284, comp_A9995_876, comp_A9_859, comp_A9992_129, comp_A3_102, comp_A3_79, comp_A9993_585, comp_A3_124, comp_A91_239, comp_A93_116, comp_A9_811, comp_A3_757, comp_A99991_336, comp_A98_66, comp_A99995_631, comp_A999_732, comp_A9996_244, comp_A995_167, comp_A98_171, comp_A3_981, comp_A9_827, comp_A9992_357, comp_A4_739, comp_A2_876, comp_A99996_412, comp_A9996_202, comp_A9993_525, comp_A7_666, comp_A92_519, comp_A99994_745, comp_A998_448, comp_A9997_490, comp_A9996_448, comp_A997_332, comp_A4_495, comp_A94_29, comp_A7_919, comp_A99997_247, comp_A993_764, comp_A9991_914, comp_A96_609, comp_A9999_832, comp_A99998_189, comp_A996_296, comp_A99999_409, comp_A99994_713, comp_A993_839, comp_A99997_833, comp_A5_327, comp_A2_894, comp_A3_587, comp_A93_629, comp_A999991_302, comp_A99997_824, comp_A9_155, comp_A5_170, comp_A97_991, comp_A995_114, comp_A5_586, comp_A98_162, comp_A991_728, comp_A9996_782, comp_A99992_505, comp_A9995_733, comp_A9991_1016, comp_A9_152, comp_A5_126, comp_A999992_426, comp_A9_784, comp_A999992_487, comp_A92_504, comp_A9994_769, comp_A95_435, comp_A999992_569, comp_A1_652, comp_A991_268, comp_A99997_799, comp_A992_599, comp_A99991_539, comp_A98_147, comp_A7_591, comp_A997_589, comp_A97_124, comp_A996_225, comp_A97_121, comp_A99995_671, comp_A9998_723, comp_A999993_9, comp_A996_92, comp_A996_222, comp_A9999_756, comp_A95_203, comp_A997_838, comp_A5_478, comp_A99997_254, comp_A99991_618, comp_A91_963, comp_A9994_288, comp_A9991_935, comp_A99997_931, comp_A98_151, comp_A4_486, comp_A3_232, comp_A9995_839, comp_A7_592, comp_A3_286, comp_A99999_486, comp_A9991_932, comp_A996_372, comp_A9_156, comp_A7_804, comp_A6_255, comp_A99991_344, comp_A8_757, comp_A993_555, comp_A999994_442, comp_A99992_671, comp_A991_479, comp_A97_610, comp_A999991_570, comp_A9_816, comp_A3_80, comp_A8_822, comp_A998_424, comp_A999993_8, comp_A9992_421, comp_A99999_549, comp_A9993_307, comp_A9996_562, comp_A996_271, comp_A992_400, comp_A94_31, comp_A99_8, comp_A3_54, comp_A2_872, comp_A92_972, comp_A3_272, comp_A999995_1015, comp_A7_605, comp_A9993_295, comp_A991_531, comp_A993_317, comp_A991_869, comp_A94_50, comp_A99994_178, comp_A8_786, comp_A3_407, comp_A6_722, comp_A99999_735, comp_A92_259, comp_A999996_390, comp_A2_901, comp_A992_675, comp_A9_821, comp_A92_503, comp_A8_536, comp_A2_124, comp_A92_250, comp_A95_497, comp_A6_406, comp_A9991_948, comp_A9999_819, comp_A3_535, comp_A998_805, comp_A92_995, comp_A9996_600, comp_A6_606, comp_A996_353, comp_A99994_600, comp_A99991_286, comp_A996_340, comp_A998_414, comp_A996_331, comp_A994_640, comp_A999_714, comp_A3_233, comp_A9_805, comp_A8_540, comp_A99996_575, comp_A993_982, comp_A9993_530, comp_A994_475, comp_A996_332, comp_A4_484, comp_A98_325, comp_A993_659, comp_A2_602, comp_A92_505, comp_A99999_58, comp_A9992_123, comp_A999992_527, comp_A9996_758, comp_A997_428, comp_A3_515, comp_A992_389, comp_A93_513, comp_A99999_558, comp_A9992_429, comp_A993_440, comp_A99996_766, comp_A999991_485, comp_A9991_1009, comp_A99999_594, comp_A993_492, comp_A96_754, comp_A993_321, comp_A999_712, comp_A997_421, comp_A9999_805, comp_A995_343, comp_A9996_570, comp_A5_653, comp_A4_445, comp_A99995_511, comp_A99991_185, comp_A99999_517, comp_A8_334, comp_A9996_737, comp_A9_845, comp_A997_339, comp_A997_243, comp_A993_683, comp_A994_543, comp_A99_13, comp_A2_22, comp_A96_818, comp_A3_350, comp_A992_528, comp_A96_271, comp_A994_365, comp_A999991_372, comp_A99999_168, comp_A95_430, comp_A8_398, comp_A994_484, comp_A999997_1009, comp_A3_415, comp_A97_174, comp_A997_549, comp_A999996_427, comp_A3_381, comp_A997_496, comp_A995_61, comp_A99_15, comp_A99_18, comp_A992_721, comp_A6_474, comp_A95_345, comp_A2_860, comp_A9_853, comp_A93_136, comp_A991_746, comp_A2_320, comp_A97_182, comp_A91_383, comp_A6_485, comp_A99995_471, comp_A93_516, comp_A99992_501, comp_A2_920, comp_A9991_961, comp_A999996_360, comp_A996_350, comp_A991_868, comp_A992_266, comp_A95_312, comp_A96_171, comp_A98_61, comp_A9994_693, comp_A994_378, comp_A99991_182, comp_A8_718, comp_A3_428, comp_A99996_862, comp_A9993_327, comp_A995_537, comp_A9_832, comp_A6_442, comp_A999996_428, comp_A94_58, comp_A997_521, comp_A996_360, comp_A99992_503, comp_A999994_457, comp_A99992_710, comp_A99991_366, comp_A993_286, comp_A999_567, comp_A99996_858, comp_A5_316, comp_A995_299, comp_A991_852, comp_A94_49, comp_A9992_105, comp_A92_247, comp_A98_68, comp_A99995_519, comp_A92_989, comp_A3_285, comp_A94_42, comp_A97_400, comp_A3_209, comp_A8_381, comp_A99_19, comp_A999997_1011, comp_A92_815, comp_A94_33, comp_A9991_937, comp_A998_499, comp_A1_554, comp_A999994_662, comp_A5_562, comp_A9997_669, comp_A997_477, comp_A9991_973, comp_A9999_248, comp_A996_245, comp_A98_1019, comp_A3_112, comp_A994_355, comp_A993_548, comp_A9991_817, comp_A92_246, comp_A3_27, comp_A8_810, comp_A99994_682, comp_A993_612, comp_A9992_99, comp_A9996_610, comp_A997_620, comp_A994_477, comp_A9999_293, comp_A8_404, comp_A996_318, comp_A95_274, comp_A1_601, comp_A92_562, comp_A99997_252, comp_A9996_694, comp_A3_305, comp_A997_334, comp_A999994_507, comp_A99993_647, comp_A992_308, comp_A99992_810, comp_A9993_652, comp_A997_403, comp_A93_651, comp_A999991_306, comp_A991_720, comp_A9992_107, comp_A9_851, comp_A9992_103, comp_A2_869, comp_A997_578, comp_A998_302, comp_A99991_660, comp_A6_644, comp_A2_285, comp_A995_202, comp_A8_818, comp_A999995_1012, comp_A997_956, comp_A999992_388, comp_A93_687, comp_A999995_1008, comp_A996_292, comp_A991_250, comp_A95_354, comp_A9994_711, comp_A9994_295, comp_A5_505, comp_A94_35, comp_A999994_547, comp_A9993_685, comp_A93_718, comp_A9991_956, comp_A993_484, comp_A1_708, comp_A9991_990, comp_A3_283, comp_A998_641, comp_A92_377, comp_A99994_383, comp_A999992_484, comp_A9_160, comp_A997_422, comp_A2_862, comp_A96_180, comp_A99997_843, comp_A9994_704, comp_A98_240, comp_A3_992, comp_A9994_881, comp_A2_827, comp_A999997_1012, comp_A994_549, comp_A97_171, comp_A9993_313, comp_A4_545, comp_A996_200, comp_A3_247, comp_A995_185, comp_A998_559, comp_A9999_767, comp_A99996_551, comp_A6_701, comp_A992_817, comp_A93_115, comp_A9991_962, comp_A99993_596, comp_A93_98, comp_A99994_807, comp_A96_264, comp_A92_500, comp_A9996_693, comp_A99993_630, comp_A99996_513, comp_A997_451, comp_A9992_161, comp_A2_114, comp_A995_493, comp_A99996_188, comp_A3_116, comp_A99996_839, comp_A2_9, comp_A93_544, comp_A3_812, comp_A997_373, comp_A99999_423, comp_A9991_955, comp_A9998_906, comp_A999996_461, comp_A999_585, comp_A5_753, comp_A99993_51, comp_A92_255, comp_A7_856, comp_A9_829, comp_A99995_559, comp_A2_33, comp_A99999_545, comp_A9992_436, comp_A997_666, comp_A94_37, comp_A9991_1011, comp_A99991_408, comp_A996_343, comp_A9999_560, comp_A996_263, comp_A9996_763, comp_A99992_660, comp_A1_642, comp_A9999_419, comp_A7_643, comp_A99992_736, comp_A9_61, comp_A6_394, comp_A99999_406, comp_A3_565, comp_A997_381, comp_A99992_538, comp_A99994_755, comp_A8_484, comp_A99992_655, comp_A991_451, comp_A99995_531, comp_A3_386, comp_A9998_389, comp_A994_390, comp_A97_201, comp_A3_750, comp_A995_34, comp_A994_677, comp_A93_720, comp_A99997_149, comp_A3_588, comp_A98_120, comp_A9_151, comp_A996_244, comp_A9999_786, comp_A99992_744, comp_A97_968, comp_A9993_626, comp_A99998_187, comp_A99994_612, comp_A9991_982, comp_A2_918, comp_A996_304, comp_A99_5, comp_A9991_693, comp_A99_21, comp_A9991_931, comp_A3_103, comp_A998_676, comp_A9_486, comp_A92_528, comp_A7_460, comp_A999994_411, comp_A93_722, comp_A98_153, comp_A996_231, comp_A999_516, comp_A991_373, comp_A9993_658, comp_A999992_474, comp_A999995_1014, comp_A9995_441, comp_A996_327, comp_A1_684, comp_A99999_443, comp_A9996_623, comp_A9_150, comp_A997_713, comp_A9991_965, comp_A999992_432, comp_A999996_726, comp_A993_258, comp_A8_335, comp_A999_656, comp_A991_735, comp_A996_203, comp_A93_546, comp_A99996_508, comp_A99996_263, comp_A9996_431, comp_A96_22, comp_A94_30, comp_A999_711, comp_A9_840, comp_A91_210, comp_A9997_587, comp_A2_713, comp_A999996_685, comp_A2_844, comp_A997_399, comp_A9993_561, comp_A991_391, comp_A6_286, comp_A99992_711, comp_A9991_921, comp_A3_55, comp_A9_157, comp_A8_657, comp_A99994_586, comp_A991_797, comp_A997_394, comp_A96_766, comp_A9993_581, comp_A9998_661, comp_A99993_699, comp_A9996_707, comp_A99997_955, comp_A991_647, comp_A996_185, comp_A999992_536, comp_A93_92, comp_A1_581, comp_A991_486, comp_A993_621, comp_A999992_339, comp_A7_767, comp_A99993_85, comp_A92_574, comp_A3_867, comp_A98_270, comp_A93_119, comp_A992_234, comp_A92_992, comp_A991_644, comp_A3_662, comp_A996_311, comp_A994_457, comp_A9993_539, comp_A99997_946, comp_A997_299, comp_A99992_670, comp_A94_32, comp_A1_741, comp_A994_524, comp_A9997_340, comp_A997_696, comp_A99994_727, comp_A994_644, comp_A996_369, comp_A9991_995, comp_A5_492, comp_A998_230, comp_A93_532, comp_A999_337, comp_A95_388, comp_A3_127, comp_A6_452, comp_A4_332, comp_A999996_581, comp_A8_875, comp_A97_207, comp_A9993_671, comp_A9999_59, comp_A991_777, comp_A9991_699, or_0, or_1, or_2, or_3, or_4, or_5, or_6, or_7, or_8, or_9, or_10, or_11, or_12, or_13, or_14, or_15, or_16, or_17, or_18, or_19, or_20, or_21, or_22, or_23, or_24
);

input [0:0] comp_A1_649;
input [0:0] comp_A2_29;
input [0:0] comp_A3_322;
input [0:0] comp_A4_504;
input [0:0] comp_A5_495;
input [0:0] comp_A6_624;
input [0:0] comp_A7_593;
input [0:0] comp_A1_220;
input [0:0] comp_A4_472;
input [0:0] comp_A8_701;
input [0:0] comp_A9_178;
input [0:0] comp_A91_362;
input [0:0] comp_A92_263;
input [0:0] comp_A93_529;
input [0:0] comp_A94_40;
input [0:0] comp_A7_795;
input [0:0] comp_A95_118;
input [0:0] comp_A3_541;
input [0:0] comp_A8_90;
input [0:0] comp_A96_11;
input [0:0] comp_A97_193;
input [0:0] comp_A98_202;
input [0:0] comp_A99_14;
input [0:0] comp_A2_830;
input [0:0] comp_A991_288;
input [0:0] comp_A992_452;
input [0:0] comp_A95_373;
input [0:0] comp_A8_777;
input [0:0] comp_A93_537;
input [0:0] comp_A99_11;
input [0:0] comp_A95_383;
input [0:0] comp_A993_454;
input [0:0] comp_A992_774;
input [0:0] comp_A994_302;
input [0:0] comp_A995_87;
input [0:0] comp_A98_143;
input [0:0] comp_A996_348;
input [0:0] comp_A997_750;
input [0:0] comp_A1_884;
input [0:0] comp_A997_360;
input [0:0] comp_A998_765;
input [0:0] comp_A8_726;
input [0:0] comp_A999_643;
input [0:0] comp_A3_526;
input [0:0] comp_A7_455;
input [0:0] comp_A9991_920;
input [0:0] comp_A3_300;
input [0:0] comp_A92_262;
input [0:0] comp_A9992_183;
input [0:0] comp_A991_737;
input [0:0] comp_A97_140;
input [0:0] comp_A9991_923;
input [0:0] comp_A96_873;
input [0:0] comp_A9993_513;
input [0:0] comp_A4_515;
input [0:0] comp_A9994_577;
input [0:0] comp_A94_46;
input [0:0] comp_A7_341;
input [0:0] comp_A3_687;
input [0:0] comp_A9995_483;
input [0:0] comp_A9996_660;
input [0:0] comp_A9997_526;
input [0:0] comp_A9991_943;
input [0:0] comp_A7_561;
input [0:0] comp_A993_276;
input [0:0] comp_A9998_478;
input [0:0] comp_A92_975;
input [0:0] comp_A1_727;
input [0:0] comp_A7_583;
input [0:0] comp_A995_79;
input [0:0] comp_A97_173;
input [0:0] comp_A993_665;
input [0:0] comp_A9999_801;
input [0:0] comp_A3_536;
input [0:0] comp_A999_620;
input [0:0] comp_A994_700;
input [0:0] comp_A99991_242;
input [0:0] comp_A994_712;
input [0:0] comp_A99992_806;
input [0:0] comp_A9997_570;
input [0:0] comp_A99993_119;
input [0:0] comp_A6_670;
input [0:0] comp_A994_338;
input [0:0] comp_A6_635;
input [0:0] comp_A9994_627;
input [0:0] comp_A1_881;
input [0:0] comp_A4_490;
input [0:0] comp_A92_264;
input [0:0] comp_A2_839;
input [0:0] comp_A991_760;
input [0:0] comp_A993_680;
input [0:0] comp_A99994_810;
input [0:0] comp_A98_974;
input [0:0] comp_A4_350;
input [0:0] comp_A1_738;
input [0:0] comp_A997_319;
input [0:0] comp_A7_411;
input [0:0] comp_A4_400;
input [0:0] comp_A9992_93;
input [0:0] comp_A99994_781;
input [0:0] comp_A93_726;
input [0:0] comp_A9998_769;
input [0:0] comp_A7_415;
input [0:0] comp_A9991_972;
input [0:0] comp_A993_608;
input [0:0] comp_A3_284;
input [0:0] comp_A9995_876;
input [0:0] comp_A9_859;
input [0:0] comp_A9992_129;
input [0:0] comp_A3_102;
input [0:0] comp_A3_79;
input [0:0] comp_A9993_585;
input [0:0] comp_A3_124;
input [0:0] comp_A91_239;
input [0:0] comp_A93_116;
input [0:0] comp_A9_811;
input [0:0] comp_A3_757;
input [0:0] comp_A99991_336;
input [0:0] comp_A98_66;
input [0:0] comp_A99995_631;
input [0:0] comp_A999_732;
input [0:0] comp_A9996_244;
input [0:0] comp_A995_167;
input [0:0] comp_A98_171;
input [0:0] comp_A3_981;
input [0:0] comp_A9_827;
input [0:0] comp_A9992_357;
input [0:0] comp_A4_739;
input [0:0] comp_A2_876;
input [0:0] comp_A99996_412;
input [0:0] comp_A9996_202;
input [0:0] comp_A9993_525;
input [0:0] comp_A7_666;
input [0:0] comp_A92_519;
input [0:0] comp_A99994_745;
input [0:0] comp_A998_448;
input [0:0] comp_A9997_490;
input [0:0] comp_A9996_448;
input [0:0] comp_A997_332;
input [0:0] comp_A4_495;
input [0:0] comp_A94_29;
input [0:0] comp_A7_919;
input [0:0] comp_A99997_247;
input [0:0] comp_A993_764;
input [0:0] comp_A9991_914;
input [0:0] comp_A96_609;
input [0:0] comp_A9999_832;
input [0:0] comp_A99998_189;
input [0:0] comp_A996_296;
input [0:0] comp_A99999_409;
input [0:0] comp_A99994_713;
input [0:0] comp_A993_839;
input [0:0] comp_A99997_833;
input [0:0] comp_A5_327;
input [0:0] comp_A2_894;
input [0:0] comp_A3_587;
input [0:0] comp_A93_629;
input [0:0] comp_A999991_302;
input [0:0] comp_A99997_824;
input [0:0] comp_A9_155;
input [0:0] comp_A5_170;
input [0:0] comp_A97_991;
input [0:0] comp_A995_114;
input [0:0] comp_A5_586;
input [0:0] comp_A98_162;
input [0:0] comp_A991_728;
input [0:0] comp_A9996_782;
input [0:0] comp_A99992_505;
input [0:0] comp_A9995_733;
input [0:0] comp_A9991_1016;
input [0:0] comp_A9_152;
input [0:0] comp_A5_126;
input [0:0] comp_A999992_426;
input [0:0] comp_A9_784;
input [0:0] comp_A999992_487;
input [0:0] comp_A92_504;
input [0:0] comp_A9994_769;
input [0:0] comp_A95_435;
input [0:0] comp_A999992_569;
input [0:0] comp_A1_652;
input [0:0] comp_A991_268;
input [0:0] comp_A99997_799;
input [0:0] comp_A992_599;
input [0:0] comp_A99991_539;
input [0:0] comp_A98_147;
input [0:0] comp_A7_591;
input [0:0] comp_A997_589;
input [0:0] comp_A97_124;
input [0:0] comp_A996_225;
input [0:0] comp_A97_121;
input [0:0] comp_A99995_671;
input [0:0] comp_A9998_723;
input [0:0] comp_A999993_9;
input [0:0] comp_A996_92;
input [0:0] comp_A996_222;
input [0:0] comp_A9999_756;
input [0:0] comp_A95_203;
input [0:0] comp_A997_838;
input [0:0] comp_A5_478;
input [0:0] comp_A99997_254;
input [0:0] comp_A99991_618;
input [0:0] comp_A91_963;
input [0:0] comp_A9994_288;
input [0:0] comp_A9991_935;
input [0:0] comp_A99997_931;
input [0:0] comp_A98_151;
input [0:0] comp_A4_486;
input [0:0] comp_A3_232;
input [0:0] comp_A9995_839;
input [0:0] comp_A7_592;
input [0:0] comp_A3_286;
input [0:0] comp_A99999_486;
input [0:0] comp_A9991_932;
input [0:0] comp_A996_372;
input [0:0] comp_A9_156;
input [0:0] comp_A7_804;
input [0:0] comp_A6_255;
input [0:0] comp_A99991_344;
input [0:0] comp_A8_757;
input [0:0] comp_A993_555;
input [0:0] comp_A999994_442;
input [0:0] comp_A99992_671;
input [0:0] comp_A991_479;
input [0:0] comp_A97_610;
input [0:0] comp_A999991_570;
input [0:0] comp_A9_816;
input [0:0] comp_A3_80;
input [0:0] comp_A8_822;
input [0:0] comp_A998_424;
input [0:0] comp_A999993_8;
input [0:0] comp_A9992_421;
input [0:0] comp_A99999_549;
input [0:0] comp_A9993_307;
input [0:0] comp_A9996_562;
input [0:0] comp_A996_271;
input [0:0] comp_A992_400;
input [0:0] comp_A94_31;
input [0:0] comp_A99_8;
input [0:0] comp_A3_54;
input [0:0] comp_A2_872;
input [0:0] comp_A92_972;
input [0:0] comp_A3_272;
input [0:0] comp_A999995_1015;
input [0:0] comp_A7_605;
input [0:0] comp_A9993_295;
input [0:0] comp_A991_531;
input [0:0] comp_A993_317;
input [0:0] comp_A991_869;
input [0:0] comp_A94_50;
input [0:0] comp_A99994_178;
input [0:0] comp_A8_786;
input [0:0] comp_A3_407;
input [0:0] comp_A6_722;
input [0:0] comp_A99999_735;
input [0:0] comp_A92_259;
input [0:0] comp_A999996_390;
input [0:0] comp_A2_901;
input [0:0] comp_A992_675;
input [0:0] comp_A9_821;
input [0:0] comp_A92_503;
input [0:0] comp_A8_536;
input [0:0] comp_A2_124;
input [0:0] comp_A92_250;
input [0:0] comp_A95_497;
input [0:0] comp_A6_406;
input [0:0] comp_A9991_948;
input [0:0] comp_A9999_819;
input [0:0] comp_A3_535;
input [0:0] comp_A998_805;
input [0:0] comp_A92_995;
input [0:0] comp_A9996_600;
input [0:0] comp_A6_606;
input [0:0] comp_A996_353;
input [0:0] comp_A99994_600;
input [0:0] comp_A99991_286;
input [0:0] comp_A996_340;
input [0:0] comp_A998_414;
input [0:0] comp_A996_331;
input [0:0] comp_A994_640;
input [0:0] comp_A999_714;
input [0:0] comp_A3_233;
input [0:0] comp_A9_805;
input [0:0] comp_A8_540;
input [0:0] comp_A99996_575;
input [0:0] comp_A993_982;
input [0:0] comp_A9993_530;
input [0:0] comp_A994_475;
input [0:0] comp_A996_332;
input [0:0] comp_A4_484;
input [0:0] comp_A98_325;
input [0:0] comp_A993_659;
input [0:0] comp_A2_602;
input [0:0] comp_A92_505;
input [0:0] comp_A99999_58;
input [0:0] comp_A9992_123;
input [0:0] comp_A999992_527;
input [0:0] comp_A9996_758;
input [0:0] comp_A997_428;
input [0:0] comp_A3_515;
input [0:0] comp_A992_389;
input [0:0] comp_A93_513;
input [0:0] comp_A99999_558;
input [0:0] comp_A9992_429;
input [0:0] comp_A993_440;
input [0:0] comp_A99996_766;
input [0:0] comp_A999991_485;
input [0:0] comp_A9991_1009;
input [0:0] comp_A99999_594;
input [0:0] comp_A993_492;
input [0:0] comp_A96_754;
input [0:0] comp_A993_321;
input [0:0] comp_A999_712;
input [0:0] comp_A997_421;
input [0:0] comp_A9999_805;
input [0:0] comp_A995_343;
input [0:0] comp_A9996_570;
input [0:0] comp_A5_653;
input [0:0] comp_A4_445;
input [0:0] comp_A99995_511;
input [0:0] comp_A99991_185;
input [0:0] comp_A99999_517;
input [0:0] comp_A8_334;
input [0:0] comp_A9996_737;
input [0:0] comp_A9_845;
input [0:0] comp_A997_339;
input [0:0] comp_A997_243;
input [0:0] comp_A993_683;
input [0:0] comp_A994_543;
input [0:0] comp_A99_13;
input [0:0] comp_A2_22;
input [0:0] comp_A96_818;
input [0:0] comp_A3_350;
input [0:0] comp_A992_528;
input [0:0] comp_A96_271;
input [0:0] comp_A994_365;
input [0:0] comp_A999991_372;
input [0:0] comp_A99999_168;
input [0:0] comp_A95_430;
input [0:0] comp_A8_398;
input [0:0] comp_A994_484;
input [0:0] comp_A999997_1009;
input [0:0] comp_A3_415;
input [0:0] comp_A97_174;
input [0:0] comp_A997_549;
input [0:0] comp_A999996_427;
input [0:0] comp_A3_381;
input [0:0] comp_A997_496;
input [0:0] comp_A995_61;
input [0:0] comp_A99_15;
input [0:0] comp_A99_18;
input [0:0] comp_A992_721;
input [0:0] comp_A6_474;
input [0:0] comp_A95_345;
input [0:0] comp_A2_860;
input [0:0] comp_A9_853;
input [0:0] comp_A93_136;
input [0:0] comp_A991_746;
input [0:0] comp_A2_320;
input [0:0] comp_A97_182;
input [0:0] comp_A91_383;
input [0:0] comp_A6_485;
input [0:0] comp_A99995_471;
input [0:0] comp_A93_516;
input [0:0] comp_A99992_501;
input [0:0] comp_A2_920;
input [0:0] comp_A9991_961;
input [0:0] comp_A999996_360;
input [0:0] comp_A996_350;
input [0:0] comp_A991_868;
input [0:0] comp_A992_266;
input [0:0] comp_A95_312;
input [0:0] comp_A96_171;
input [0:0] comp_A98_61;
input [0:0] comp_A9994_693;
input [0:0] comp_A994_378;
input [0:0] comp_A99991_182;
input [0:0] comp_A8_718;
input [0:0] comp_A3_428;
input [0:0] comp_A99996_862;
input [0:0] comp_A9993_327;
input [0:0] comp_A995_537;
input [0:0] comp_A9_832;
input [0:0] comp_A6_442;
input [0:0] comp_A999996_428;
input [0:0] comp_A94_58;
input [0:0] comp_A997_521;
input [0:0] comp_A996_360;
input [0:0] comp_A99992_503;
input [0:0] comp_A999994_457;
input [0:0] comp_A99992_710;
input [0:0] comp_A99991_366;
input [0:0] comp_A993_286;
input [0:0] comp_A999_567;
input [0:0] comp_A99996_858;
input [0:0] comp_A5_316;
input [0:0] comp_A995_299;
input [0:0] comp_A991_852;
input [0:0] comp_A94_49;
input [0:0] comp_A9992_105;
input [0:0] comp_A92_247;
input [0:0] comp_A98_68;
input [0:0] comp_A99995_519;
input [0:0] comp_A92_989;
input [0:0] comp_A3_285;
input [0:0] comp_A94_42;
input [0:0] comp_A97_400;
input [0:0] comp_A3_209;
input [0:0] comp_A8_381;
input [0:0] comp_A99_19;
input [0:0] comp_A999997_1011;
input [0:0] comp_A92_815;
input [0:0] comp_A94_33;
input [0:0] comp_A9991_937;
input [0:0] comp_A998_499;
input [0:0] comp_A1_554;
input [0:0] comp_A999994_662;
input [0:0] comp_A5_562;
input [0:0] comp_A9997_669;
input [0:0] comp_A997_477;
input [0:0] comp_A9991_973;
input [0:0] comp_A9999_248;
input [0:0] comp_A996_245;
input [0:0] comp_A98_1019;
input [0:0] comp_A3_112;
input [0:0] comp_A994_355;
input [0:0] comp_A993_548;
input [0:0] comp_A9991_817;
input [0:0] comp_A92_246;
input [0:0] comp_A3_27;
input [0:0] comp_A8_810;
input [0:0] comp_A99994_682;
input [0:0] comp_A993_612;
input [0:0] comp_A9992_99;
input [0:0] comp_A9996_610;
input [0:0] comp_A997_620;
input [0:0] comp_A994_477;
input [0:0] comp_A9999_293;
input [0:0] comp_A8_404;
input [0:0] comp_A996_318;
input [0:0] comp_A95_274;
input [0:0] comp_A1_601;
input [0:0] comp_A92_562;
input [0:0] comp_A99997_252;
input [0:0] comp_A9996_694;
input [0:0] comp_A3_305;
input [0:0] comp_A997_334;
input [0:0] comp_A999994_507;
input [0:0] comp_A99993_647;
input [0:0] comp_A992_308;
input [0:0] comp_A99992_810;
input [0:0] comp_A9993_652;
input [0:0] comp_A997_403;
input [0:0] comp_A93_651;
input [0:0] comp_A999991_306;
input [0:0] comp_A991_720;
input [0:0] comp_A9992_107;
input [0:0] comp_A9_851;
input [0:0] comp_A9992_103;
input [0:0] comp_A2_869;
input [0:0] comp_A997_578;
input [0:0] comp_A998_302;
input [0:0] comp_A99991_660;
input [0:0] comp_A6_644;
input [0:0] comp_A2_285;
input [0:0] comp_A995_202;
input [0:0] comp_A8_818;
input [0:0] comp_A999995_1012;
input [0:0] comp_A997_956;
input [0:0] comp_A999992_388;
input [0:0] comp_A93_687;
input [0:0] comp_A999995_1008;
input [0:0] comp_A996_292;
input [0:0] comp_A991_250;
input [0:0] comp_A95_354;
input [0:0] comp_A9994_711;
input [0:0] comp_A9994_295;
input [0:0] comp_A5_505;
input [0:0] comp_A94_35;
input [0:0] comp_A999994_547;
input [0:0] comp_A9993_685;
input [0:0] comp_A93_718;
input [0:0] comp_A9991_956;
input [0:0] comp_A993_484;
input [0:0] comp_A1_708;
input [0:0] comp_A9991_990;
input [0:0] comp_A3_283;
input [0:0] comp_A998_641;
input [0:0] comp_A92_377;
input [0:0] comp_A99994_383;
input [0:0] comp_A999992_484;
input [0:0] comp_A9_160;
input [0:0] comp_A997_422;
input [0:0] comp_A2_862;
input [0:0] comp_A96_180;
input [0:0] comp_A99997_843;
input [0:0] comp_A9994_704;
input [0:0] comp_A98_240;
input [0:0] comp_A3_992;
input [0:0] comp_A9994_881;
input [0:0] comp_A2_827;
input [0:0] comp_A999997_1012;
input [0:0] comp_A994_549;
input [0:0] comp_A97_171;
input [0:0] comp_A9993_313;
input [0:0] comp_A4_545;
input [0:0] comp_A996_200;
input [0:0] comp_A3_247;
input [0:0] comp_A995_185;
input [0:0] comp_A998_559;
input [0:0] comp_A9999_767;
input [0:0] comp_A99996_551;
input [0:0] comp_A6_701;
input [0:0] comp_A992_817;
input [0:0] comp_A93_115;
input [0:0] comp_A9991_962;
input [0:0] comp_A99993_596;
input [0:0] comp_A93_98;
input [0:0] comp_A99994_807;
input [0:0] comp_A96_264;
input [0:0] comp_A92_500;
input [0:0] comp_A9996_693;
input [0:0] comp_A99993_630;
input [0:0] comp_A99996_513;
input [0:0] comp_A997_451;
input [0:0] comp_A9992_161;
input [0:0] comp_A2_114;
input [0:0] comp_A995_493;
input [0:0] comp_A99996_188;
input [0:0] comp_A3_116;
input [0:0] comp_A99996_839;
input [0:0] comp_A2_9;
input [0:0] comp_A93_544;
input [0:0] comp_A3_812;
input [0:0] comp_A997_373;
input [0:0] comp_A99999_423;
input [0:0] comp_A9991_955;
input [0:0] comp_A9998_906;
input [0:0] comp_A999996_461;
input [0:0] comp_A999_585;
input [0:0] comp_A5_753;
input [0:0] comp_A99993_51;
input [0:0] comp_A92_255;
input [0:0] comp_A7_856;
input [0:0] comp_A9_829;
input [0:0] comp_A99995_559;
input [0:0] comp_A2_33;
input [0:0] comp_A99999_545;
input [0:0] comp_A9992_436;
input [0:0] comp_A997_666;
input [0:0] comp_A94_37;
input [0:0] comp_A9991_1011;
input [0:0] comp_A99991_408;
input [0:0] comp_A996_343;
input [0:0] comp_A9999_560;
input [0:0] comp_A996_263;
input [0:0] comp_A9996_763;
input [0:0] comp_A99992_660;
input [0:0] comp_A1_642;
input [0:0] comp_A9999_419;
input [0:0] comp_A7_643;
input [0:0] comp_A99992_736;
input [0:0] comp_A9_61;
input [0:0] comp_A6_394;
input [0:0] comp_A99999_406;
input [0:0] comp_A3_565;
input [0:0] comp_A997_381;
input [0:0] comp_A99992_538;
input [0:0] comp_A99994_755;
input [0:0] comp_A8_484;
input [0:0] comp_A99992_655;
input [0:0] comp_A991_451;
input [0:0] comp_A99995_531;
input [0:0] comp_A3_386;
input [0:0] comp_A9998_389;
input [0:0] comp_A994_390;
input [0:0] comp_A97_201;
input [0:0] comp_A3_750;
input [0:0] comp_A995_34;
input [0:0] comp_A994_677;
input [0:0] comp_A93_720;
input [0:0] comp_A99997_149;
input [0:0] comp_A3_588;
input [0:0] comp_A98_120;
input [0:0] comp_A9_151;
input [0:0] comp_A996_244;
input [0:0] comp_A9999_786;
input [0:0] comp_A99992_744;
input [0:0] comp_A97_968;
input [0:0] comp_A9993_626;
input [0:0] comp_A99998_187;
input [0:0] comp_A99994_612;
input [0:0] comp_A9991_982;
input [0:0] comp_A2_918;
input [0:0] comp_A996_304;
input [0:0] comp_A99_5;
input [0:0] comp_A9991_693;
input [0:0] comp_A99_21;
input [0:0] comp_A9991_931;
input [0:0] comp_A3_103;
input [0:0] comp_A998_676;
input [0:0] comp_A9_486;
input [0:0] comp_A92_528;
input [0:0] comp_A7_460;
input [0:0] comp_A999994_411;
input [0:0] comp_A93_722;
input [0:0] comp_A98_153;
input [0:0] comp_A996_231;
input [0:0] comp_A999_516;
input [0:0] comp_A991_373;
input [0:0] comp_A9993_658;
input [0:0] comp_A999992_474;
input [0:0] comp_A999995_1014;
input [0:0] comp_A9995_441;
input [0:0] comp_A996_327;
input [0:0] comp_A1_684;
input [0:0] comp_A99999_443;
input [0:0] comp_A9996_623;
input [0:0] comp_A9_150;
input [0:0] comp_A997_713;
input [0:0] comp_A9991_965;
input [0:0] comp_A999992_432;
input [0:0] comp_A999996_726;
input [0:0] comp_A993_258;
input [0:0] comp_A8_335;
input [0:0] comp_A999_656;
input [0:0] comp_A991_735;
input [0:0] comp_A996_203;
input [0:0] comp_A93_546;
input [0:0] comp_A99996_508;
input [0:0] comp_A99996_263;
input [0:0] comp_A9996_431;
input [0:0] comp_A96_22;
input [0:0] comp_A94_30;
input [0:0] comp_A999_711;
input [0:0] comp_A9_840;
input [0:0] comp_A91_210;
input [0:0] comp_A9997_587;
input [0:0] comp_A2_713;
input [0:0] comp_A999996_685;
input [0:0] comp_A2_844;
input [0:0] comp_A997_399;
input [0:0] comp_A9993_561;
input [0:0] comp_A991_391;
input [0:0] comp_A6_286;
input [0:0] comp_A99992_711;
input [0:0] comp_A9991_921;
input [0:0] comp_A3_55;
input [0:0] comp_A9_157;
input [0:0] comp_A8_657;
input [0:0] comp_A99994_586;
input [0:0] comp_A991_797;
input [0:0] comp_A997_394;
input [0:0] comp_A96_766;
input [0:0] comp_A9993_581;
input [0:0] comp_A9998_661;
input [0:0] comp_A99993_699;
input [0:0] comp_A9996_707;
input [0:0] comp_A99997_955;
input [0:0] comp_A991_647;
input [0:0] comp_A996_185;
input [0:0] comp_A999992_536;
input [0:0] comp_A93_92;
input [0:0] comp_A1_581;
input [0:0] comp_A991_486;
input [0:0] comp_A993_621;
input [0:0] comp_A999992_339;
input [0:0] comp_A7_767;
input [0:0] comp_A99993_85;
input [0:0] comp_A92_574;
input [0:0] comp_A3_867;
input [0:0] comp_A98_270;
input [0:0] comp_A93_119;
input [0:0] comp_A992_234;
input [0:0] comp_A92_992;
input [0:0] comp_A991_644;
input [0:0] comp_A3_662;
input [0:0] comp_A996_311;
input [0:0] comp_A994_457;
input [0:0] comp_A9993_539;
input [0:0] comp_A99997_946;
input [0:0] comp_A997_299;
input [0:0] comp_A99992_670;
input [0:0] comp_A94_32;
input [0:0] comp_A1_741;
input [0:0] comp_A994_524;
input [0:0] comp_A9997_340;
input [0:0] comp_A997_696;
input [0:0] comp_A99994_727;
input [0:0] comp_A994_644;
input [0:0] comp_A996_369;
input [0:0] comp_A9991_995;
input [0:0] comp_A5_492;
input [0:0] comp_A998_230;
input [0:0] comp_A93_532;
input [0:0] comp_A999_337;
input [0:0] comp_A95_388;
input [0:0] comp_A3_127;
input [0:0] comp_A6_452;
input [0:0] comp_A4_332;
input [0:0] comp_A999996_581;
input [0:0] comp_A8_875;
input [0:0] comp_A97_207;
input [0:0] comp_A9993_671;
input [0:0] comp_A9999_59;
input [0:0] comp_A991_777;
input [0:0] comp_A9991_699;
output [0:0] or_0;
output [0:0] or_1;
output [0:0] or_2;
output [0:0] or_3;
output [0:0] or_4;
output [0:0] or_5;
output [0:0] or_6;
output [0:0] or_7;
output [0:0] or_8;
output [0:0] or_9;
output [0:0] or_10;
output [0:0] or_11;
output [0:0] or_12;
output [0:0] or_13;
output [0:0] or_14;
output [0:0] or_15;
output [0:0] or_16;
output [0:0] or_17;
output [0:0] or_18;
output [0:0] or_19;
output [0:0] or_20;
output [0:0] or_21;
output [0:0] or_22;
output [0:0] or_23;
output [0:0] or_24;

wire [0:0] and_0;
wire [0:0] and_1;
wire [0:0] and_2;
wire [0:0] and_3;
wire [0:0] and_4;
wire [0:0] and_5;
wire [0:0] and_6;
wire [0:0] and_7;
wire [0:0] and_8;
wire [0:0] and_9;
wire [0:0] and_10;
wire [0:0] and_11;
wire [0:0] and_12;
wire [0:0] and_13;
wire [0:0] and_14;
wire [0:0] and_15;
wire [0:0] and_16;
wire [0:0] and_17;
wire [0:0] and_18;
wire [0:0] and_19;
wire [0:0] and_20;
wire [0:0] and_21;
wire [0:0] and_22;
wire [0:0] and_23;
wire [0:0] and_24;
wire [0:0] and_25;
wire [0:0] and_26;
wire [0:0] and_27;
wire [0:0] and_28;
wire [0:0] and_29;
wire [0:0] and_30;
wire [0:0] and_31;
wire [0:0] and_32;
wire [0:0] and_33;
wire [0:0] and_34;
wire [0:0] and_35;
wire [0:0] and_36;
wire [0:0] and_37;
wire [0:0] and_38;
wire [0:0] and_39;
wire [0:0] and_40;
wire [0:0] and_41;
wire [0:0] and_42;
wire [0:0] and_43;
wire [0:0] and_44;
wire [0:0] and_45;
wire [0:0] and_46;
wire [0:0] and_47;
wire [0:0] and_48;
wire [0:0] and_49;
wire [0:0] and_50;
wire [0:0] and_51;
wire [0:0] and_52;
wire [0:0] and_53;
wire [0:0] and_54;
wire [0:0] and_55;
wire [0:0] and_56;
wire [0:0] and_57;
wire [0:0] and_58;
wire [0:0] and_59;
wire [0:0] and_60;
wire [0:0] and_61;
wire [0:0] and_62;
wire [0:0] and_63;
wire [0:0] and_64;
wire [0:0] and_65;
wire [0:0] and_66;
wire [0:0] and_67;
wire [0:0] and_68;
wire [0:0] and_69;
wire [0:0] and_70;
wire [0:0] and_71;
wire [0:0] and_72;
wire [0:0] and_73;
wire [0:0] and_74;
wire [0:0] and_75;
wire [0:0] and_76;
wire [0:0] and_77;
wire [0:0] and_78;
wire [0:0] and_79;
wire [0:0] and_80;
wire [0:0] and_81;
wire [0:0] and_82;
wire [0:0] and_83;
wire [0:0] and_84;
wire [0:0] and_85;
wire [0:0] and_86;
wire [0:0] and_87;
wire [0:0] and_88;
wire [0:0] and_89;
wire [0:0] and_90;
wire [0:0] and_91;
wire [0:0] and_92;
wire [0:0] and_93;
wire [0:0] and_94;
wire [0:0] and_95;
wire [0:0] and_96;
wire [0:0] and_97;
wire [0:0] and_98;
wire [0:0] and_99;
wire [0:0] and_100;
wire [0:0] and_101;
wire [0:0] and_102;
wire [0:0] and_103;
wire [0:0] and_104;
wire [0:0] and_105;
wire [0:0] and_106;
wire [0:0] and_107;
wire [0:0] and_108;
wire [0:0] and_109;
wire [0:0] and_110;
wire [0:0] and_111;
wire [0:0] and_112;
wire [0:0] and_113;
wire [0:0] and_114;
wire [0:0] and_115;
wire [0:0] and_116;
wire [0:0] and_117;
wire [0:0] and_118;
wire [0:0] and_119;
wire [0:0] and_120;
wire [0:0] and_121;
wire [0:0] and_122;
wire [0:0] and_123;
wire [0:0] and_124;
wire [0:0] and_125;
wire [0:0] and_126;
wire [0:0] and_127;
wire [0:0] and_128;
wire [0:0] and_129;
wire [0:0] and_130;
wire [0:0] and_131;
wire [0:0] and_132;
wire [0:0] and_133;
wire [0:0] and_134;
wire [0:0] and_135;
wire [0:0] and_136;
wire [0:0] and_137;
wire [0:0] and_138;
wire [0:0] and_139;
wire [0:0] and_140;
wire [0:0] and_141;
wire [0:0] and_142;
wire [0:0] and_143;
wire [0:0] and_144;
wire [0:0] and_145;
wire [0:0] and_146;
wire [0:0] and_147;
wire [0:0] and_148;
wire [0:0] and_149;
wire [0:0] and_150;
wire [0:0] and_151;
wire [0:0] and_152;
wire [0:0] and_153;
wire [0:0] and_154;
wire [0:0] and_155;
wire [0:0] and_156;
wire [0:0] and_157;
wire [0:0] and_158;
wire [0:0] and_159;
wire [0:0] and_160;
wire [0:0] and_161;
wire [0:0] and_162;
wire [0:0] and_163;
wire [0:0] and_164;
wire [0:0] and_165;
wire [0:0] and_166;
wire [0:0] and_167;
wire [0:0] and_168;
wire [0:0] and_169;
wire [0:0] and_170;
wire [0:0] and_171;
wire [0:0] and_172;
wire [0:0] and_173;
wire [0:0] and_174;
wire [0:0] and_175;
wire [0:0] and_176;
wire [0:0] and_177;
wire [0:0] and_178;
wire [0:0] and_179;
wire [0:0] and_180;
wire [0:0] and_181;
wire [0:0] and_182;
wire [0:0] and_183;
wire [0:0] and_184;
wire [0:0] and_185;
wire [0:0] and_186;
wire [0:0] and_187;
wire [0:0] and_188;
wire [0:0] and_189;
wire [0:0] and_190;
wire [0:0] and_191;
wire [0:0] and_192;
wire [0:0] and_193;
wire [0:0] and_194;
wire [0:0] and_195;
wire [0:0] and_196;
wire [0:0] and_197;
wire [0:0] and_198;
wire [0:0] and_199;
wire [0:0] and_200;
wire [0:0] and_201;
wire [0:0] and_202;
wire [0:0] and_203;
wire [0:0] and_204;
wire [0:0] and_205;
wire [0:0] and_206;
wire [0:0] and_207;
wire [0:0] and_208;
wire [0:0] and_209;
wire [0:0] and_210;
wire [0:0] and_211;
wire [0:0] and_212;
wire [0:0] and_213;
wire [0:0] and_214;
wire [0:0] and_215;
wire [0:0] and_216;
wire [0:0] and_217;
wire [0:0] and_218;
wire [0:0] and_219;
wire [0:0] and_220;
wire [0:0] and_221;
wire [0:0] and_222;
wire [0:0] and_223;
wire [0:0] and_224;
wire [0:0] and_225;
wire [0:0] and_226;
wire [0:0] and_227;
wire [0:0] and_228;
wire [0:0] and_229;
wire [0:0] and_230;
wire [0:0] and_231;
wire [0:0] and_232;
wire [0:0] and_233;
wire [0:0] and_234;
wire [0:0] and_235;
wire [0:0] and_236;
wire [0:0] and_237;
wire [0:0] and_238;
wire [0:0] and_239;
wire [0:0] and_240;
wire [0:0] and_241;
wire [0:0] and_242;
wire [0:0] and_243;
wire [0:0] and_244;
wire [0:0] and_245;
wire [0:0] and_246;
wire [0:0] and_247;
wire [0:0] and_248;
wire [0:0] and_249;
wire [0:0] and_250;
wire [0:0] and_251;
wire [0:0] and_252;
wire [0:0] and_253;
wire [0:0] and_254;
wire [0:0] and_255;
wire [0:0] and_256;
wire [0:0] and_257;
wire [0:0] and_258;
wire [0:0] and_259;
wire [0:0] and_260;
wire [0:0] and_261;
wire [0:0] and_262;
wire [0:0] and_263;
wire [0:0] and_264;
wire [0:0] and_265;
wire [0:0] and_266;
wire [0:0] and_267;
wire [0:0] and_268;
wire [0:0] and_269;
wire [0:0] and_270;
wire [0:0] and_271;
wire [0:0] and_272;
wire [0:0] and_273;
wire [0:0] and_274;
wire [0:0] and_275;
wire [0:0] and_276;
wire [0:0] and_277;
wire [0:0] and_278;
wire [0:0] and_279;
wire [0:0] and_280;
wire [0:0] and_281;
wire [0:0] and_282;
wire [0:0] and_283;
wire [0:0] and_284;
wire [0:0] and_285;
wire [0:0] and_286;
wire [0:0] and_287;
wire [0:0] and_288;
wire [0:0] and_289;
wire [0:0] and_290;
wire [0:0] and_291;
wire [0:0] and_292;
wire [0:0] and_293;
wire [0:0] and_294;
wire [0:0] and_295;
wire [0:0] and_296;
wire [0:0] and_297;
wire [0:0] and_298;
wire [0:0] and_299;
wire [0:0] and_300;
wire [0:0] and_301;
wire [0:0] and_302;
wire [0:0] and_303;
wire [0:0] and_304;
wire [0:0] and_305;
wire [0:0] and_306;
wire [0:0] and_307;
wire [0:0] and_308;
wire [0:0] and_309;
wire [0:0] and_310;
wire [0:0] and_311;
wire [0:0] and_312;
wire [0:0] and_313;
wire [0:0] and_314;
wire [0:0] and_315;
wire [0:0] and_316;
wire [0:0] and_317;
wire [0:0] and_318;
wire [0:0] and_319;
wire [0:0] and_320;
wire [0:0] and_321;
wire [0:0] and_322;
wire [0:0] and_323;
wire [0:0] and_324;
wire [0:0] and_325;
wire [0:0] and_326;
wire [0:0] and_327;
wire [0:0] and_328;
wire [0:0] and_329;
wire [0:0] and_330;
wire [0:0] and_331;
wire [0:0] and_332;
wire [0:0] and_333;
wire [0:0] and_334;
wire [0:0] and_335;
wire [0:0] and_336;
wire [0:0] and_337;
wire [0:0] and_338;
wire [0:0] and_339;
wire [0:0] and_340;
wire [0:0] and_341;
wire [0:0] and_342;
wire [0:0] and_343;
wire [0:0] and_344;
wire [0:0] and_345;
wire [0:0] and_346;
wire [0:0] and_347;
wire [0:0] and_348;
wire [0:0] and_349;
wire [0:0] and_350;
wire [0:0] and_351;
wire [0:0] and_352;
wire [0:0] and_353;
wire [0:0] and_354;
wire [0:0] and_355;
wire [0:0] and_356;
wire [0:0] and_357;
wire [0:0] and_358;
wire [0:0] and_359;
wire [0:0] and_360;
wire [0:0] and_361;
wire [0:0] and_362;
wire [0:0] and_363;
wire [0:0] and_364;
wire [0:0] and_365;
wire [0:0] and_366;
wire [0:0] and_367;
wire [0:0] and_368;
wire [0:0] and_369;
wire [0:0] and_370;
wire [0:0] and_371;
wire [0:0] and_372;
wire [0:0] and_373;
wire [0:0] and_374;
wire [0:0] and_375;
wire [0:0] and_376;
wire [0:0] and_377;
wire [0:0] and_378;
wire [0:0] and_379;
wire [0:0] and_380;
wire [0:0] and_381;
wire [0:0] and_382;
wire [0:0] and_383;
wire [0:0] and_384;
wire [0:0] and_385;
wire [0:0] and_386;
wire [0:0] and_387;
wire [0:0] and_388;
wire [0:0] and_389;
wire [0:0] and_390;
wire [0:0] and_391;
wire [0:0] and_392;
wire [0:0] and_393;
wire [0:0] and_394;
wire [0:0] and_395;
wire [0:0] and_396;
wire [0:0] and_397;
wire [0:0] and_398;
wire [0:0] and_399;
wire [0:0] and_400;
wire [0:0] and_401;
wire [0:0] and_402;
wire [0:0] and_403;
wire [0:0] and_404;
wire [0:0] and_405;
wire [0:0] and_406;
wire [0:0] and_407;
wire [0:0] and_408;
wire [0:0] and_409;
wire [0:0] and_410;
wire [0:0] and_411;
wire [0:0] and_412;
wire [0:0] and_413;
wire [0:0] and_414;
wire [0:0] and_415;
wire [0:0] and_416;
wire [0:0] and_417;
wire [0:0] and_418;
wire [0:0] and_419;
wire [0:0] and_420;
wire [0:0] and_421;
wire [0:0] and_422;
wire [0:0] and_423;
wire [0:0] and_424;
wire [0:0] and_425;
wire [0:0] and_426;
wire [0:0] and_427;
wire [0:0] and_428;
wire [0:0] and_429;
wire [0:0] and_430;
wire [0:0] and_431;
wire [0:0] and_432;
wire [0:0] and_433;
wire [0:0] and_434;
wire [0:0] and_435;
wire [0:0] and_436;
wire [0:0] and_437;
wire [0:0] and_438;
wire [0:0] and_439;
wire [0:0] and_440;
wire [0:0] and_441;
wire [0:0] and_442;
wire [0:0] and_443;
wire [0:0] and_444;
wire [0:0] and_445;
wire [0:0] and_446;
wire [0:0] and_447;
wire [0:0] and_448;
wire [0:0] and_449;
wire [0:0] and_450;
wire [0:0] and_451;
wire [0:0] and_452;
wire [0:0] and_453;
wire [0:0] and_454;
wire [0:0] and_455;
wire [0:0] and_456;
wire [0:0] and_457;
wire [0:0] and_458;
wire [0:0] and_459;
wire [0:0] and_460;
wire [0:0] and_461;
wire [0:0] and_462;
wire [0:0] and_463;
wire [0:0] and_464;
wire [0:0] and_465;
wire [0:0] and_466;
wire [0:0] and_467;
wire [0:0] and_468;
wire [0:0] and_469;
wire [0:0] and_470;
wire [0:0] and_471;
wire [0:0] and_472;
wire [0:0] and_473;
wire [0:0] and_474;
wire [0:0] and_475;
wire [0:0] and_476;
wire [0:0] and_477;
wire [0:0] and_478;
wire [0:0] and_479;
wire [0:0] and_480;
wire [0:0] and_481;
wire [0:0] and_482;
wire [0:0] and_483;
wire [0:0] and_484;
wire [0:0] and_485;
wire [0:0] and_486;
wire [0:0] and_487;
wire [0:0] and_488;
wire [0:0] and_489;
wire [0:0] and_490;
wire [0:0] and_491;
wire [0:0] and_492;
wire [0:0] and_493;
wire [0:0] and_494;
wire [0:0] and_495;
wire [0:0] and_496;
wire [0:0] and_497;
wire [0:0] and_498;
wire [0:0] and_499;
wire [0:0] and_500;
wire [0:0] and_501;
wire [0:0] and_502;
wire [0:0] and_503;
wire [0:0] and_504;
wire [0:0] and_505;
wire [0:0] and_506;
wire [0:0] and_507;
wire [0:0] and_508;
wire [0:0] and_509;
wire [0:0] and_510;
wire [0:0] and_511;
wire [0:0] and_512;
wire [0:0] and_513;
wire [0:0] and_514;
wire [0:0] and_515;
wire [0:0] and_516;
wire [0:0] and_517;
wire [0:0] and_518;
wire [0:0] and_519;
wire [0:0] and_520;
wire [0:0] and_521;
wire [0:0] and_522;
wire [0:0] and_523;
wire [0:0] and_524;
wire [0:0] and_525;
wire [0:0] and_526;
wire [0:0] and_527;
wire [0:0] and_528;
wire [0:0] and_529;
wire [0:0] and_530;
wire [0:0] and_531;
wire [0:0] and_532;
wire [0:0] and_533;
wire [0:0] and_534;
wire [0:0] and_535;
wire [0:0] and_536;
wire [0:0] and_537;
wire [0:0] and_538;
wire [0:0] and_539;
wire [0:0] and_540;
wire [0:0] and_541;
wire [0:0] and_542;
wire [0:0] and_543;
wire [0:0] and_544;
wire [0:0] and_545;
wire [0:0] and_546;
wire [0:0] and_547;
wire [0:0] and_548;
wire [0:0] and_549;
wire [0:0] and_550;
wire [0:0] and_551;
wire [0:0] and_552;
wire [0:0] and_553;
wire [0:0] and_554;
wire [0:0] and_555;
wire [0:0] and_556;
wire [0:0] and_557;
wire [0:0] and_558;
wire [0:0] and_559;
wire [0:0] and_560;
wire [0:0] and_561;
wire [0:0] and_562;
wire [0:0] and_563;
wire [0:0] and_564;
wire [0:0] and_565;
wire [0:0] and_566;
wire [0:0] and_567;
wire [0:0] and_568;
wire [0:0] and_569;
wire [0:0] and_570;
wire [0:0] and_571;
wire [0:0] and_572;
wire [0:0] and_573;
wire [0:0] and_574;
wire [0:0] and_575;
wire [0:0] and_576;
wire [0:0] and_577;
wire [0:0] and_578;
wire [0:0] and_579;
wire [0:0] and_580;
wire [0:0] and_581;
wire [0:0] and_582;
wire [0:0] and_583;
wire [0:0] and_584;
wire [0:0] and_585;
wire [0:0] and_586;
wire [0:0] and_587;
wire [0:0] and_588;
wire [0:0] and_589;
wire [0:0] and_590;
wire [0:0] and_591;
wire [0:0] and_592;
wire [0:0] and_593;
wire [0:0] and_594;
wire [0:0] and_595;
wire [0:0] and_596;
wire [0:0] and_597;
wire [0:0] and_598;
wire [0:0] and_599;
wire [0:0] and_600;
wire [0:0] and_601;
wire [0:0] and_602;
wire [0:0] and_603;
wire [0:0] and_604;
wire [0:0] and_605;
wire [0:0] and_606;
wire [0:0] and_607;
wire [0:0] and_608;
wire [0:0] and_609;
wire [0:0] and_610;
wire [0:0] and_611;
wire [0:0] and_612;
wire [0:0] and_613;
wire [0:0] and_614;
wire [0:0] and_615;
wire [0:0] and_616;
wire [0:0] and_617;
wire [0:0] and_618;
wire [0:0] and_619;
wire [0:0] and_620;
wire [0:0] and_621;
wire [0:0] and_622;
wire [0:0] and_623;
wire [0:0] and_624;
wire [0:0] and_625;
wire [0:0] and_626;
wire [0:0] and_627;
wire [0:0] and_628;
wire [0:0] and_629;
wire [0:0] and_630;
wire [0:0] and_631;
wire [0:0] and_632;
wire [0:0] and_633;
wire [0:0] and_634;
wire [0:0] and_635;
wire [0:0] and_636;
wire [0:0] and_637;
wire [0:0] and_638;
wire [0:0] and_639;
wire [0:0] and_640;
wire [0:0] and_641;
wire [0:0] and_642;
wire [0:0] and_643;
wire [0:0] and_644;
wire [0:0] and_645;
wire [0:0] and_646;
wire [0:0] and_647;
wire [0:0] and_648;
wire [0:0] and_649;
wire [0:0] and_650;
wire [0:0] and_651;
wire [0:0] and_652;
wire [0:0] and_653;
wire [0:0] and_654;
wire [0:0] and_655;
wire [0:0] and_656;
wire [0:0] and_657;
wire [0:0] and_658;
wire [0:0] and_659;
wire [0:0] and_660;
wire [0:0] and_661;
wire [0:0] and_662;
wire [0:0] and_663;
wire [0:0] and_664;
wire [0:0] and_665;
wire [0:0] and_666;
wire [0:0] and_667;
wire [0:0] and_668;
wire [0:0] and_669;
wire [0:0] and_670;
wire [0:0] and_671;
wire [0:0] and_672;
wire [0:0] and_673;
wire [0:0] and_674;
wire [0:0] and_675;
wire [0:0] and_676;
wire [0:0] and_677;
wire [0:0] and_678;
wire [0:0] and_679;
wire [0:0] and_680;
wire [0:0] and_681;
wire [0:0] and_682;
wire [0:0] and_683;
wire [0:0] and_684;
wire [0:0] and_685;
wire [0:0] and_686;
wire [0:0] and_687;
wire [0:0] and_688;
wire [0:0] and_689;
wire [0:0] and_690;
wire [0:0] and_691;
wire [0:0] and_692;
wire [0:0] and_693;
wire [0:0] and_694;
wire [0:0] and_695;
wire [0:0] and_696;
wire [0:0] and_697;
wire [0:0] and_698;
wire [0:0] and_699;
wire [0:0] and_700;
wire [0:0] and_701;
wire [0:0] and_702;
wire [0:0] and_703;
wire [0:0] and_704;
wire [0:0] and_705;
wire [0:0] and_706;
wire [0:0] and_707;
wire [0:0] and_708;
wire [0:0] and_709;
wire [0:0] and_710;
wire [0:0] and_711;
wire [0:0] and_712;
wire [0:0] and_713;
wire [0:0] and_714;
wire [0:0] and_715;
wire [0:0] and_716;
wire [0:0] and_717;
wire [0:0] and_718;
wire [0:0] and_719;
wire [0:0] and_720;
wire [0:0] and_721;
wire [0:0] and_722;
wire [0:0] and_723;
wire [0:0] and_724;
wire [0:0] and_725;
wire [0:0] and_726;
wire [0:0] and_727;
wire [0:0] and_728;
wire [0:0] and_729;
wire [0:0] and_730;
wire [0:0] and_731;
wire [0:0] and_732;
wire [0:0] and_733;
wire [0:0] and_734;
wire [0:0] and_735;
wire [0:0] and_736;
wire [0:0] and_737;
wire [0:0] and_738;
wire [0:0] and_739;
wire [0:0] and_740;
wire [0:0] and_741;
wire [0:0] and_742;
wire [0:0] and_743;
wire [0:0] and_744;
wire [0:0] and_745;
wire [0:0] and_746;
wire [0:0] and_747;
wire [0:0] and_748;
wire [0:0] and_749;
wire [0:0] and_750;
wire [0:0] and_751;
wire [0:0] and_752;
wire [0:0] and_753;
wire [0:0] and_754;
wire [0:0] and_755;
wire [0:0] and_756;
wire [0:0] and_757;
wire [0:0] and_758;
wire [0:0] and_759;

assign and_0 = comp_A1_649 & comp_A2_29 & comp_A3_322 & ~(comp_A4_504) & ~(comp_A5_495) & ~(comp_A6_624);

assign and_1 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & ~(comp_A9_178) & comp_A7_795 & ~(comp_A95_118) & comp_A8_90;

assign and_2 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & ~(comp_A4_350) & ~(comp_A4_400) & ~(comp_A9998_769);

assign and_3 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & comp_A93_537 & comp_A9995_876 & comp_A9_859 & ~(comp_A9992_129);

assign and_4 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & ~(comp_A93_537) & comp_A3_102 & comp_A3_79 & ~(comp_A9993_585);

assign and_5 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & comp_A93_116 & comp_A9_811 & ~(comp_A3_757);

assign and_6 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & comp_A9996_244 & comp_A995_167 & ~(comp_A98_171);

assign and_7 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & ~(comp_A9996_244) & comp_A9_827 & comp_A9992_357;

assign and_8 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A9_811 & comp_A2_876 & comp_A99996_412 & ~(comp_A9996_202) & ~(comp_A7_666);

assign and_9 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A9_811) & comp_A2_876 & comp_A99996_412 & comp_A92_519 & comp_A99994_745;

assign and_10 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & comp_A998_448 & comp_A9997_490 & ~(comp_A9996_448);

assign and_11 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & ~(comp_A998_448) & comp_A4_495 & ~(comp_A94_29);

assign and_12 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & ~(comp_A998_448) & ~(comp_A4_495) & comp_A7_919;

assign and_13 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & comp_A99999_409 & comp_A99994_713 & ~(comp_A993_839);

assign and_14 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & ~(comp_A99999_409) & comp_A5_327 & comp_A2_894;

assign and_15 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & comp_A9996_782 & comp_A99992_505 & ~(comp_A9995_733);

assign and_16 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & ~(comp_A991_288) & comp_A95_383 & comp_A993_454;

assign and_17 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & ~(comp_A991_288) & comp_A95_383 & ~(comp_A994_302);

assign and_18 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & ~(comp_A991_288) & ~(comp_A95_383) & comp_A995_87 & comp_A98_143;

assign and_19 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & comp_A1_884 & comp_A997_360 & ~(comp_A998_765);

assign and_20 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & ~(comp_A1_884) & comp_A999_643 & comp_A3_526;

assign and_21 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & ~(comp_A997_750) & ~(comp_A9991_920) & ~(comp_A9992_183);

assign and_22 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & comp_A97_140 & ~(comp_A9991_923) & comp_A4_515 & comp_A9994_577;

assign and_23 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & ~(comp_A97_140) & comp_A94_46 & ~(comp_A7_341) & ~(comp_A9995_483);

assign and_24 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & comp_A9991_943 & comp_A7_561 & comp_A993_276;

assign and_25 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & comp_A995_79 & comp_A97_173 & comp_A993_665;

assign and_26 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & ~(comp_A995_79) & comp_A3_536 & comp_A999_620;

assign and_27 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & comp_A994_712 & comp_A99992_806 & ~(comp_A9997_570) & ~(comp_A994_338) & ~(comp_A6_635);

assign and_28 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & comp_A2_839 & comp_A991_760 & comp_A993_680;

assign and_29 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & comp_A2_839 & ~(comp_A991_760) & comp_A99994_810;

assign and_30 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & comp_A2_839 & ~(comp_A991_760) & ~(comp_A98_974);

assign or_0 = and_0 | and_1 | and_2 | and_3 | and_4 | and_5 | and_6 | and_7 | and_8 | and_9 | and_10 | and_11 | and_12 | and_13 | and_14 | and_15 | and_16 | and_17 | and_18 | and_19 | and_20 | and_21 | and_22 | and_23 | and_24 | and_25 | and_26 | and_27 | and_28 | and_29 | and_30;

assign and_31 = comp_A1_649 & comp_A2_29 & comp_A3_322 & ~(comp_A4_504) & comp_A5_495;

assign and_32 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & comp_A9_178 & comp_A91_362 & comp_A92_263 & comp_A93_529 & comp_A94_40;

assign and_33 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & ~(comp_A4_350) & comp_A4_400 & comp_A9992_93 & ~(comp_A99994_781);

assign and_34 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & ~(comp_A4_350) & comp_A4_400 & ~(comp_A9992_93) & ~(comp_A93_726);

assign and_35 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & ~(comp_A4_350) & ~(comp_A4_400) & comp_A9998_769 & ~(comp_A7_415);

assign and_36 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & ~(comp_A93_537) & comp_A3_102 & ~(comp_A3_79);

assign and_37 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & comp_A93_116 & comp_A9_811 & comp_A3_757 & comp_A99991_336;

assign and_38 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & comp_A93_116 & ~(comp_A9_811) & comp_A99995_631;

assign and_39 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & comp_A9996_244 & ~(comp_A995_167) & ~(comp_A3_981);

assign and_40 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A9_811 & comp_A2_876 & comp_A99996_412 & comp_A9996_202 & comp_A9993_525;

assign and_41 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A9_811) & comp_A2_876 & comp_A99996_412 & comp_A92_519 & ~(comp_A99994_745);

assign and_42 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & comp_A998_448 & ~(comp_A9997_490) & comp_A997_332;

assign and_43 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & ~(comp_A998_448) & comp_A4_495 & comp_A94_29;

assign and_44 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & comp_A99997_247 & comp_A993_764 & comp_A9991_914 & ~(comp_A96_609);

assign and_45 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & comp_A99997_247 & comp_A993_764 & ~(comp_A9991_914) & comp_A9999_832;

assign and_46 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & comp_A99997_247 & ~(comp_A993_764) & ~(comp_A99998_189);

assign and_47 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & comp_A99997_247 & ~(comp_A993_764) & comp_A996_296;

assign and_48 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A9_811 & comp_A93_629 & ~(comp_A999991_302) & comp_A995_114 & comp_A5_586 & ~(comp_A98_162);

assign and_49 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & comp_A999991_302 & comp_A99997_824 & comp_A9_155 & comp_A5_170;

assign and_50 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & comp_A999991_302 & comp_A99997_824 & ~(comp_A9_155) & comp_A97_991;

assign and_51 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & comp_A995_114 & ~(comp_A5_586) & comp_A991_728;

assign and_52 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & comp_A9996_782 & ~(comp_A99992_505) & ~(comp_A9991_1016);

assign and_53 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & ~(comp_A9996_782) & comp_A9_152 & comp_A5_126;

assign and_54 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & ~(comp_A9996_782) & ~(comp_A9_152) & ~(comp_A999992_426);

assign and_55 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & ~(comp_A995_114) & ~(comp_A9_784);

assign and_56 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & comp_A9_784 & comp_A999992_487 & comp_A92_504;

assign and_57 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & comp_A991_288 & comp_A992_452 & ~(comp_A95_373) & ~(comp_A8_777);

assign and_58 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & comp_A991_288 & ~(comp_A992_452) & comp_A93_537 & comp_A99_11;

assign and_59 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & ~(comp_A991_288) & ~(comp_A95_383) & comp_A995_87 & ~(comp_A98_143);

assign and_60 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & comp_A1_884 & comp_A997_360 & comp_A998_765;

assign and_61 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & comp_A1_884 & ~(comp_A997_360) & comp_A8_726;

assign and_62 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & ~(comp_A1_884) & ~(comp_A999_643) & ~(comp_A7_455);

assign and_63 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & ~(comp_A997_750) & comp_A9991_920 & comp_A3_300;

assign and_64 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & comp_A97_140 & ~(comp_A9991_923) & comp_A4_515 & ~(comp_A9994_577);

assign and_65 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & ~(comp_A97_140) & comp_A94_46 & comp_A7_341 & ~(comp_A3_687);

assign and_66 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & ~(comp_A97_140) & ~(comp_A94_46) & ~(comp_A9996_660) & comp_A9997_526;

assign and_67 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & comp_A9991_943 & ~(comp_A7_561) & ~(comp_A92_975) & comp_A7_583;

assign and_68 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & comp_A995_79 & ~(comp_A97_173) & ~(comp_A9999_801);

assign and_69 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & ~(comp_A995_79) & comp_A3_536 & ~(comp_A999_620);

assign and_70 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & comp_A994_712 & ~(comp_A99992_806);

assign and_71 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & comp_A994_712 & ~(comp_A9997_570) & ~(comp_A994_338) & comp_A6_635;

assign and_72 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & ~(comp_A994_712) & comp_A9994_627 & comp_A1_881;

assign and_73 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & ~(comp_A994_712) & comp_A9994_627 & ~(comp_A4_490) & comp_A92_264;

assign and_74 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & comp_A2_839 & comp_A991_760 & ~(comp_A993_680);

assign and_75 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & comp_A2_839 & ~(comp_A991_760) & ~(comp_A99994_810) & comp_A98_974;

assign and_76 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & comp_A4_350 & comp_A1_738 & comp_A997_319;

assign and_77 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & comp_A4_350 & ~(comp_A1_738) & ~(comp_A7_411);

assign or_1 = and_31 | and_32 | and_33 | and_34 | and_35 | and_36 | and_37 | and_38 | and_39 | and_40 | and_41 | and_42 | and_43 | and_44 | and_45 | and_46 | and_47 | and_48 | and_49 | and_50 | and_51 | and_52 | and_53 | and_54 | and_55 | and_56 | and_57 | and_58 | and_59 | and_60 | and_61 | and_62 | and_63 | and_64 | and_65 | and_66 | and_67 | and_68 | and_69 | and_70 | and_71 | and_72 | and_73 | and_74 | and_75 | and_76 | and_77;

assign and_78 = comp_A1_649 & comp_A2_29 & comp_A3_322 & ~(comp_A4_504) & ~(comp_A5_495) & comp_A6_624;

assign and_79 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & comp_A9_178 & comp_A91_362 & comp_A92_263 & comp_A93_529 & ~(comp_A94_40);

assign and_80 = comp_A1_649 & ~(comp_A2_29) & comp_A1_220 & ~(comp_A4_472) & comp_A8_701;

assign and_81 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & ~(comp_A4_350) & comp_A4_400 & comp_A9992_93 & comp_A99994_781;

assign and_82 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & ~(comp_A4_350) & comp_A4_400 & ~(comp_A9992_93) & comp_A93_726;

assign and_83 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & ~(comp_A93_537) & ~(comp_A3_102) & comp_A3_124;

assign and_84 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & comp_A9996_244 & comp_A995_167 & comp_A98_171;

assign and_85 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & ~(comp_A9996_244) & ~(comp_A9_827) & ~(comp_A4_739);

assign and_86 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A9_811 & comp_A2_876 & comp_A99996_412 & comp_A9996_202 & ~(comp_A9993_525);

assign and_87 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & comp_A99999_409 & ~(comp_A99994_713) & ~(comp_A99997_833);

assign and_88 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & ~(comp_A99999_409) & ~(comp_A5_327) & comp_A3_587;

assign and_89 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & comp_A995_114 & ~(comp_A5_586) & ~(comp_A991_728);

assign and_90 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & comp_A991_288 & comp_A992_452 & comp_A95_373;

assign and_91 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & comp_A991_288 & comp_A992_452 & comp_A8_777;

assign and_92 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & comp_A991_288 & ~(comp_A992_452) & comp_A93_537 & ~(comp_A99_11);

assign and_93 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & ~(comp_A991_288) & comp_A95_383 & ~(comp_A993_454) & comp_A994_302;

assign and_94 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & ~(comp_A991_288) & ~(comp_A95_383) & ~(comp_A995_87) & comp_A996_348;

assign and_95 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & comp_A1_884 & ~(comp_A997_360) & ~(comp_A8_726);

assign and_96 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & ~(comp_A1_884) & comp_A999_643 & ~(comp_A3_526);

assign and_97 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & comp_A997_750 & ~(comp_A1_884) & ~(comp_A999_643) & comp_A7_455;

assign and_98 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & ~(comp_A997_750) & comp_A9991_920 & ~(comp_A3_300) & comp_A92_262;

assign and_99 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & comp_A97_140 & comp_A9991_923 & comp_A96_873 & comp_A9993_513;

assign and_100 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & comp_A97_140 & ~(comp_A9991_923) & ~(comp_A4_515);

assign and_101 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & ~(comp_A97_140) & comp_A94_46 & comp_A7_341 & comp_A3_687;

assign and_102 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & ~(comp_A97_140) & comp_A94_46 & ~(comp_A7_341) & comp_A9995_483;

assign and_103 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & comp_A9991_943 & comp_A7_561 & ~(comp_A993_276) & ~(comp_A9998_478);

assign and_104 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & comp_A9991_943 & ~(comp_A7_561) & comp_A92_975 & ~(comp_A1_727);

assign and_105 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & ~(comp_A995_79) & ~(comp_A3_536) & comp_A994_700;

assign and_106 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & comp_A994_712 & comp_A99992_806 & ~(comp_A9997_570) & comp_A994_338;

assign and_107 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & ~(comp_A994_712) & comp_A9994_627 & ~(comp_A1_881) & comp_A4_490;

assign and_108 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & comp_A4_350 & comp_A1_738 & ~(comp_A997_319);

assign and_109 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & comp_A4_350 & ~(comp_A1_738) & comp_A7_411;

assign or_2 = and_78 | and_79 | and_80 | and_81 | and_82 | and_83 | and_84 | and_85 | and_86 | and_87 | and_88 | and_89 | and_90 | and_91 | and_92 | and_93 | and_94 | and_95 | and_96 | and_97 | and_98 | and_99 | and_100 | and_101 | and_102 | and_103 | and_104 | and_105 | and_106 | and_107 | and_108 | and_109;

assign and_110 = comp_A1_649 & comp_A2_29 & ~(comp_A3_322) & ~(comp_A7_593);

assign and_111 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & comp_A9_178 & comp_A91_362 & ~(comp_A92_263);

assign and_112 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & ~(comp_A9_178) & ~(comp_A7_795);

assign and_113 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & ~(comp_A9_178) & comp_A95_118 & ~(comp_A3_541);

assign and_114 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & ~(comp_A9_178) & ~(comp_A95_118) & ~(comp_A8_90) & comp_A96_11;

assign and_115 = comp_A1_649 & ~(comp_A2_29) & comp_A1_220 & ~(comp_A4_472) & ~(comp_A8_701);

assign and_116 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & ~(comp_A93_537) & ~(comp_A3_102) & ~(comp_A3_124) & comp_A91_239;

assign and_117 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & comp_A93_116 & comp_A9_811 & comp_A3_757 & ~(comp_A99991_336);

assign and_118 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & comp_A93_116 & ~(comp_A9_811) & ~(comp_A99995_631) & comp_A999_732;

assign and_119 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & ~(comp_A9996_244) & comp_A9_827 & ~(comp_A9992_357);

assign and_120 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A9_811 & comp_A2_876 & comp_A99996_412 & ~(comp_A9996_202) & comp_A7_666;

assign and_121 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & comp_A99997_247 & comp_A993_764 & ~(comp_A9991_914) & ~(comp_A9999_832);

assign and_122 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & comp_A99999_409 & comp_A99994_713 & comp_A993_839;

assign and_123 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & comp_A99999_409 & ~(comp_A99994_713) & comp_A99997_833;

assign and_124 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A9_811 & comp_A93_629 & ~(comp_A999991_302) & comp_A995_114 & comp_A5_586 & comp_A98_162;

assign and_125 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & comp_A9996_782 & comp_A99992_505 & comp_A9995_733;

assign and_126 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & comp_A995_114 & ~(comp_A9_784) & comp_A999992_569;

assign and_127 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & comp_A9_784 & comp_A999992_487 & ~(comp_A92_504) & comp_A9994_769;

assign and_128 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & comp_A9_784 & ~(comp_A999992_487) & ~(comp_A95_435);

assign and_129 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & ~(comp_A97_140) & ~(comp_A94_46) & ~(comp_A9996_660) & ~(comp_A9997_526);

assign and_130 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & comp_A9991_943 & ~(comp_A7_561) & ~(comp_A92_975) & ~(comp_A7_583);

assign and_131 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & comp_A995_79 & comp_A97_173 & ~(comp_A993_665);

assign and_132 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & comp_A995_79 & ~(comp_A97_173) & comp_A9999_801;

assign and_133 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & comp_A994_712 & comp_A99992_806 & comp_A9997_570 & ~(comp_A99993_119);

assign and_134 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & comp_A994_712 & comp_A99992_806 & comp_A9997_570 & comp_A6_670;

assign or_3 = and_110 | and_111 | and_112 | and_113 | and_114 | and_115 | and_116 | and_117 | and_118 | and_119 | and_120 | and_121 | and_122 | and_123 | and_124 | and_125 | and_126 | and_127 | and_128 | and_129 | and_130 | and_131 | and_132 | and_133 | and_134;

assign and_135 = comp_A1_649 & comp_A2_29 & comp_A3_322 & comp_A4_504;

assign and_136 = comp_A1_649 & comp_A2_29 & ~(comp_A3_322) & comp_A7_593;

assign and_137 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & comp_A9_178 & ~(comp_A91_362);

assign and_138 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & comp_A9_178 & comp_A92_263 & ~(comp_A93_529);

assign and_139 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & ~(comp_A9_178) & comp_A7_795 & comp_A95_118 & comp_A3_541;

assign and_140 = comp_A1_649 & ~(comp_A2_29) & ~(comp_A1_220) & ~(comp_A9_178) & comp_A7_795 & ~(comp_A95_118) & ~(comp_A8_90) & ~(comp_A96_11);

assign and_141 = comp_A1_649 & ~(comp_A2_29) & comp_A1_220 & comp_A4_472;

assign and_142 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & ~(comp_A99991_242) & ~(comp_A2_839) & ~(comp_A4_350) & ~(comp_A4_400) & comp_A9998_769 & comp_A7_415;

assign and_143 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & comp_A93_537 & ~(comp_A9995_876);

assign and_144 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & comp_A93_537 & ~(comp_A9_859);

assign and_145 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & comp_A93_537 & comp_A9992_129;

assign and_146 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & ~(comp_A93_537) & comp_A3_102 & comp_A3_79 & comp_A9993_585;

assign and_147 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & comp_A3_284 & ~(comp_A93_537) & ~(comp_A3_102) & ~(comp_A3_124) & ~(comp_A91_239);

assign and_148 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & comp_A93_116 & ~(comp_A9_811) & ~(comp_A99995_631) & ~(comp_A999_732);

assign and_149 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & comp_A9996_244 & ~(comp_A995_167) & comp_A3_981;

assign and_150 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & comp_A993_608 & ~(comp_A3_284) & ~(comp_A93_116) & ~(comp_A9996_244) & ~(comp_A9_827) & comp_A4_739;

assign and_151 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A9_811) & comp_A2_876 & comp_A99996_412 & ~(comp_A92_519);

assign and_152 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & comp_A998_448 & comp_A9997_490 & comp_A9996_448;

assign and_153 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & comp_A998_448 & ~(comp_A9997_490) & ~(comp_A997_332);

assign and_154 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & comp_A2_876 & ~(comp_A99996_412) & ~(comp_A998_448) & ~(comp_A4_495) & ~(comp_A7_919);

assign and_155 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & comp_A99997_247 & comp_A993_764 & comp_A9991_914 & comp_A96_609;

assign and_156 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & comp_A99997_247 & ~(comp_A993_764) & comp_A99998_189 & ~(comp_A996_296);

assign and_157 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & ~(comp_A99999_409) & comp_A5_327 & ~(comp_A2_894);

assign and_158 = ~(comp_A1_649) & ~(comp_A97_193) & comp_A9991_972 & ~(comp_A993_608) & ~(comp_A2_876) & ~(comp_A99997_247) & ~(comp_A99999_409) & ~(comp_A5_327) & ~(comp_A3_587);

assign and_159 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A9_811) & comp_A93_629 & ~(comp_A999991_302) & comp_A995_114 & comp_A5_586;

assign and_160 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & comp_A999991_302 & ~(comp_A99997_824);

assign and_161 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & comp_A999991_302 & comp_A9_155 & ~(comp_A5_170);

assign and_162 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & comp_A999991_302 & ~(comp_A9_155) & ~(comp_A97_991);

assign and_163 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & comp_A9996_782 & ~(comp_A99992_505) & comp_A9991_1016;

assign and_164 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & ~(comp_A9996_782) & comp_A9_152 & ~(comp_A5_126);

assign and_165 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & comp_A93_629 & ~(comp_A999991_302) & ~(comp_A995_114) & ~(comp_A9996_782) & ~(comp_A9_152) & comp_A999992_426;

assign and_166 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & comp_A995_114 & ~(comp_A9_784) & ~(comp_A999992_569);

assign and_167 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & comp_A9_784 & comp_A999992_487 & ~(comp_A92_504) & ~(comp_A9994_769);

assign and_168 = ~(comp_A1_649) & ~(comp_A97_193) & ~(comp_A9991_972) & ~(comp_A93_629) & comp_A9_784 & ~(comp_A999992_487) & comp_A95_435;

assign and_169 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & comp_A991_288 & ~(comp_A992_452) & ~(comp_A93_537);

assign and_170 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & comp_A2_830 & ~(comp_A991_288) & ~(comp_A95_383) & ~(comp_A995_87) & ~(comp_A996_348);

assign and_171 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & ~(comp_A997_750) & comp_A9991_920 & ~(comp_A3_300) & ~(comp_A92_262);

assign and_172 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & comp_A99_14 & ~(comp_A2_830) & ~(comp_A997_750) & ~(comp_A9991_920) & comp_A9992_183;

assign and_173 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & comp_A97_140 & comp_A9991_923 & ~(comp_A96_873);

assign and_174 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & comp_A97_140 & comp_A9991_923 & ~(comp_A9993_513);

assign and_175 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & comp_A991_737 & ~(comp_A97_140) & ~(comp_A94_46) & comp_A9996_660;

assign and_176 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & comp_A9991_943 & comp_A7_561 & ~(comp_A993_276) & comp_A9998_478;

assign and_177 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & comp_A9991_943 & ~(comp_A7_561) & comp_A92_975 & comp_A1_727;

assign and_178 = ~(comp_A1_649) & comp_A97_193 & comp_A98_202 & ~(comp_A99_14) & ~(comp_A991_737) & ~(comp_A9991_943) & ~(comp_A995_79) & ~(comp_A3_536) & ~(comp_A994_700);

assign and_179 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & comp_A994_712 & comp_A99992_806 & comp_A9997_570 & comp_A99993_119 & ~(comp_A6_670);

assign and_180 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & ~(comp_A994_712) & ~(comp_A9994_627);

assign and_181 = ~(comp_A1_649) & comp_A97_193 & ~(comp_A98_202) & comp_A99991_242 & ~(comp_A994_712) & ~(comp_A1_881) & ~(comp_A4_490) & ~(comp_A92_264);

assign or_4 = and_135 | and_136 | and_137 | and_138 | and_139 | and_140 | and_141 | and_142 | and_143 | and_144 | and_145 | and_146 | and_147 | and_148 | and_149 | and_150 | and_151 | and_152 | and_153 | and_154 | and_155 | and_156 | and_157 | and_158 | and_159 | and_160 | and_161 | and_162 | and_163 | and_164 | and_165 | and_166 | and_167 | and_168 | and_169 | and_170 | and_171 | and_172 | and_173 | and_174 | and_175 | and_176 | and_177 | and_178 | and_179 | and_180 | and_181;

assign and_182 = comp_A2_29 & comp_A92_263 & comp_A9991_972 & comp_A1_652 & ~(comp_A991_268) & ~(comp_A99991_539) & ~(comp_A98_147);

assign and_183 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & comp_A97_124 & ~(comp_A996_225);

assign and_184 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & ~(comp_A97_124) & comp_A99995_671 & ~(comp_A9998_723) & ~(comp_A999993_9);

assign and_185 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & ~(comp_A996_222) & ~(comp_A91_963) & ~(comp_A9994_288);

assign and_186 = comp_A997_360 & comp_A9991_972 & ~(comp_A98_66) & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & comp_A4_486 & ~(comp_A3_232);

assign and_187 = comp_A9991_972 & comp_A2_876 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & ~(comp_A991_869) & ~(comp_A99999_735);

assign and_188 = comp_A9991_972 & comp_A9993_525 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & comp_A92_972 & comp_A3_272;

assign and_189 = comp_A9991_972 & comp_A995_114 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & comp_A92_995 & comp_A9996_600;

assign and_190 = comp_A9991_972 & comp_A995_114 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & comp_A92_995 & ~(comp_A6_606);

assign and_191 = comp_A9991_972 & ~(comp_A995_114) & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & comp_A92_995 & ~(comp_A996_353) & comp_A99991_286;

assign and_192 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & comp_A3_286 & comp_A99999_486 & ~(comp_A9991_932);

assign and_193 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & comp_A3_286 & ~(comp_A99999_486) & comp_A996_372;

assign and_194 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & comp_A99991_344 & comp_A8_757 & comp_A993_555;

assign and_195 = ~(comp_A9992_93) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & ~(comp_A99991_344) & comp_A97_610 & ~(comp_A9_816);

assign and_196 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & ~(comp_A99991_344) & ~(comp_A97_610) & comp_A3_80;

assign and_197 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & comp_A998_424 & comp_A999993_8 & ~(comp_A9992_421);

assign and_198 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & comp_A998_424 & comp_A999993_8 & comp_A99999_549;

assign and_199 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & comp_A998_424 & comp_A999993_8 & ~(comp_A9993_307);

assign and_200 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & comp_A9996_562 & comp_A996_271 & comp_A992_400 & comp_A94_31;

assign and_201 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & comp_A9996_562 & comp_A996_271 & ~(comp_A992_400) & ~(comp_A99_8);

assign and_202 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & ~(comp_A92_972) & comp_A7_605 & ~(comp_A9993_295);

assign and_203 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & ~(comp_A92_972) & ~(comp_A7_605) & comp_A991_531;

assign and_204 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & comp_A991_869 & comp_A94_50 & ~(comp_A99994_178) & comp_A8_786;

assign and_205 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & comp_A991_869 & comp_A94_50 & ~(comp_A99994_178) & comp_A3_407;

assign and_206 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & comp_A991_869 & ~(comp_A94_50) & ~(comp_A6_722);

assign and_207 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & ~(comp_A991_869) & comp_A99999_735 & comp_A92_259;

assign and_208 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & comp_A992_675 & comp_A9_821 & comp_A92_503;

assign and_209 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & ~(comp_A992_675) & comp_A2_124 & ~(comp_A92_250);

assign and_210 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & ~(comp_A992_675) & ~(comp_A2_124) & comp_A95_497;

assign and_211 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & ~(comp_A2_901) & ~(comp_A6_406) & comp_A3_535 & comp_A998_805;

assign and_212 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & ~(comp_A92_995) & comp_A996_340 & ~(comp_A998_414) & ~(comp_A996_331);

assign and_213 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & ~(comp_A92_995) & ~(comp_A996_340) & comp_A994_640;

assign and_214 = ~(comp_A93_537) & ~(comp_A9991_972) & comp_A92_503 & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & comp_A997_421 & ~(comp_A9999_805) & ~(comp_A995_343);

assign and_215 = comp_A93_537 & ~(comp_A9991_972) & ~(comp_A3_233) & ~(comp_A9993_530) & ~(comp_A99999_594) & ~(comp_A993_321);

assign and_216 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & comp_A9996_758 & comp_A997_428 & comp_A3_515 & comp_A992_389;

assign or_5 = and_182 | and_183 | and_184 | and_185 | and_186 | and_187 | and_188 | and_189 | and_190 | and_191 | and_192 | and_193 | and_194 | and_195 | and_196 | and_197 | and_198 | and_199 | and_200 | and_201 | and_202 | and_203 | and_204 | and_205 | and_206 | and_207 | and_208 | and_209 | and_210 | and_211 | and_212 | and_213 | and_214 | and_215 | and_216;

assign and_217 = comp_A2_29 & comp_A92_263 & comp_A9991_972 & comp_A1_652 & comp_A991_268 & comp_A99997_799;

assign and_218 = comp_A2_29 & comp_A92_263 & comp_A9991_972 & comp_A1_652 & comp_A991_268 & ~(comp_A992_599);

assign and_219 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & ~(comp_A9999_756) & comp_A997_838 & ~(comp_A5_478) & comp_A99997_254;

assign and_220 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & ~(comp_A9999_756) & ~(comp_A997_838) & comp_A99991_618;

assign and_221 = ~(comp_A92_263) & comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & ~(comp_A2_901) & comp_A6_406 & ~(comp_A9999_819);

assign and_222 = comp_A997_360 & comp_A9991_972 & comp_A98_66 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & comp_A4_486 & ~(comp_A3_232);

assign and_223 = comp_A9991_972 & ~(comp_A2_876) & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & ~(comp_A991_869) & ~(comp_A99999_735);

assign and_224 = comp_A9991_972 & ~(comp_A995_114) & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & comp_A92_995 & comp_A996_353 & ~(comp_A99994_600);

assign and_225 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & comp_A99991_344 & comp_A8_757 & ~(comp_A993_555) & comp_A999994_442;

assign and_226 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & comp_A99991_344 & ~(comp_A8_757) & comp_A99992_671 & comp_A991_479;

assign and_227 = comp_A9992_93 & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & ~(comp_A99991_344) & comp_A97_610 & ~(comp_A999991_570);

assign and_228 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & ~(comp_A99991_344) & ~(comp_A97_610) & ~(comp_A3_80) & ~(comp_A8_822);

assign and_229 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & ~(comp_A92_972) & ~(comp_A7_605) & ~(comp_A991_531);

assign and_230 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & comp_A991_869 & comp_A94_50 & comp_A99994_178;

assign and_231 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & comp_A991_869 & comp_A94_50 & ~(comp_A8_786) & ~(comp_A3_407);

assign and_232 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & comp_A991_869 & ~(comp_A94_50) & comp_A6_722;

assign and_233 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & comp_A993_317 & ~(comp_A991_869) & comp_A99999_735 & ~(comp_A92_259);

assign and_234 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & comp_A992_675 & ~(comp_A9_821) & ~(comp_A8_536);

assign and_235 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & ~(comp_A2_901) & ~(comp_A6_406) & comp_A3_535 & ~(comp_A998_805);

assign and_236 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & ~(comp_A92_995) & comp_A996_340 & ~(comp_A998_414) & comp_A996_331;

assign and_237 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & ~(comp_A92_995) & ~(comp_A996_340) & ~(comp_A994_640) & ~(comp_A999_714);

assign and_238 = comp_A93_537 & ~(comp_A9991_972) & comp_A99998_189 & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A99999_594 & comp_A993_492;

assign and_239 = ~(comp_A9991_972) & ~(comp_A999992_426) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & ~(comp_A9996_758) & comp_A9992_429 & ~(comp_A993_440);

assign and_240 = ~(comp_A9991_972) & comp_A9_784 & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & comp_A996_332;

assign and_241 = ~(comp_A93_537) & ~(comp_A9991_972) & comp_A92_503 & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & comp_A997_421 & comp_A9999_805;

assign and_242 = ~(comp_A93_537) & ~(comp_A9991_972) & comp_A92_503 & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & comp_A997_421 & comp_A995_343;

assign and_243 = ~(comp_A93_537) & ~(comp_A9991_972) & ~(comp_A92_503) & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & comp_A997_421 & comp_A9996_570 & ~(comp_A5_653);

assign and_244 = comp_A93_537 & ~(comp_A9991_972) & ~(comp_A3_233) & ~(comp_A9993_530) & ~(comp_A99999_594) & comp_A993_321;

assign and_245 = ~(comp_A93_537) & ~(comp_A9991_972) & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & ~(comp_A997_421) & comp_A4_445;

assign and_246 = ~(comp_A93_537) & ~(comp_A9991_972) & ~(comp_A3_233) & ~(comp_A9993_530) & ~(comp_A999_712) & ~(comp_A99995_511);

assign and_247 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & comp_A996_332 & comp_A4_484 & ~(comp_A98_325);

assign and_248 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & ~(comp_A996_332) & comp_A993_659 & comp_A2_602 & comp_A92_505 & ~(comp_A99999_58);

assign and_249 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & ~(comp_A996_332) & ~(comp_A993_659) & comp_A9992_123;

assign and_250 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & comp_A9996_758 & comp_A997_428 & ~(comp_A3_515);

assign and_251 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & comp_A9996_758 & comp_A997_428 & ~(comp_A992_389);

assign and_252 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & ~(comp_A9996_758) & ~(comp_A9992_429) & ~(comp_A999991_485) & comp_A9991_1009;

assign or_6 = and_217 | and_218 | and_219 | and_220 | and_221 | and_222 | and_223 | and_224 | and_225 | and_226 | and_227 | and_228 | and_229 | and_230 | and_231 | and_232 | and_233 | and_234 | and_235 | and_236 | and_237 | and_238 | and_239 | and_240 | and_241 | and_242 | and_243 | and_244 | and_245 | and_246 | and_247 | and_248 | and_249 | and_250 | and_251 | and_252;

assign and_253 = comp_A2_29 & comp_A92_263 & comp_A9991_972 & comp_A1_652 & comp_A991_268 & ~(comp_A99997_799) & comp_A992_599;

assign and_254 = comp_A2_29 & comp_A92_263 & comp_A9991_972 & comp_A1_652 & ~(comp_A991_268) & ~(comp_A99991_539) & comp_A98_147;

assign and_255 = ~(comp_A2_29) & comp_A8_701 & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & comp_A9999_756 & comp_A95_203;

assign and_256 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & ~(comp_A9999_756) & comp_A997_838 & ~(comp_A5_478) & ~(comp_A99997_254);

assign and_257 = comp_A92_263 & comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & ~(comp_A2_901) & comp_A6_406 & comp_A9991_948;

assign and_258 = comp_A9991_972 & comp_A9993_525 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & comp_A92_972 & ~(comp_A3_272);

assign and_259 = comp_A997_360 & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & ~(comp_A4_486) & ~(comp_A9995_839);

assign and_260 = comp_A997_360 & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & ~(comp_A4_486) & ~(comp_A7_592);

assign and_261 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & ~(comp_A3_286) & ~(comp_A9_156) & ~(comp_A6_255);

assign and_262 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & comp_A99991_344 & ~(comp_A8_757) & comp_A99992_671 & ~(comp_A991_479);

assign and_263 = ~(comp_A9992_93) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & ~(comp_A99991_344) & comp_A97_610 & comp_A9_816;

assign and_264 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & comp_A998_424 & comp_A999993_8 & comp_A9992_421 & ~(comp_A99999_549) & comp_A9993_307;

assign and_265 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & comp_A9996_562 & comp_A996_271 & comp_A992_400 & ~(comp_A94_31);

assign and_266 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & comp_A9996_562 & comp_A996_271 & ~(comp_A992_400) & comp_A99_8;

assign and_267 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & comp_A9996_562 & ~(comp_A996_271) & ~(comp_A3_54) & ~(comp_A2_872);

assign and_268 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & ~(comp_A92_972) & comp_A7_605 & comp_A9993_295;

assign and_269 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & comp_A992_675 & comp_A9_821 & ~(comp_A92_503);

assign and_270 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & ~(comp_A992_675) & ~(comp_A2_124) & ~(comp_A95_497);

assign and_271 = ~(comp_A93_537) & ~(comp_A9991_972) & ~(comp_A92_503) & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & comp_A997_421 & comp_A9996_570 & comp_A5_653;

assign and_272 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & comp_A9996_758 & ~(comp_A997_428) & ~(comp_A93_513) & ~(comp_A99999_558);

assign and_273 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & ~(comp_A9996_758) & comp_A9992_429 & comp_A993_440 & ~(comp_A99996_766);

assign or_7 = and_253 | and_254 | and_255 | and_256 | and_257 | and_258 | and_259 | and_260 | and_261 | and_262 | and_263 | and_264 | and_265 | and_266 | and_267 | and_268 | and_269 | and_270 | and_271 | and_272 | and_273;

assign and_274 = comp_A2_29 & ~(comp_A92_263) & comp_A9991_972 & comp_A1_652 & ~(comp_A7_591);

assign and_275 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & comp_A97_124 & comp_A996_225 & ~(comp_A97_121);

assign and_276 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & ~(comp_A97_124) & ~(comp_A99995_671) & comp_A996_92;

assign and_277 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & comp_A9999_756 & ~(comp_A95_203);

assign and_278 = ~(comp_A2_29) & ~(comp_A8_701) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & comp_A9999_756;

assign and_279 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & ~(comp_A9999_756) & comp_A997_838 & comp_A5_478;

assign and_280 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & comp_A996_222 & ~(comp_A9999_756) & ~(comp_A997_838) & ~(comp_A99991_618);

assign and_281 = comp_A92_263 & comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & ~(comp_A2_901) & comp_A6_406 & ~(comp_A9991_948);

assign and_282 = comp_A9991_972 & ~(comp_A9993_525) & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & comp_A92_972 & ~(comp_A999995_1015);

assign and_283 = comp_A9991_972 & comp_A995_114 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & comp_A92_995 & ~(comp_A9996_600) & comp_A6_606;

assign and_284 = comp_A9991_972 & ~(comp_A995_114) & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & comp_A92_995 & ~(comp_A996_353) & ~(comp_A99991_286);

assign and_285 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & ~(comp_A3_286) & comp_A9_156 & ~(comp_A7_804);

assign and_286 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & ~(comp_A99991_344) & ~(comp_A97_610) & ~(comp_A3_80) & comp_A8_822;

assign and_287 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & comp_A998_424 & ~(comp_A999993_8);

assign and_288 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & comp_A9996_562 & ~(comp_A996_271) & ~(comp_A3_54) & comp_A2_872;

assign and_289 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & ~(comp_A992_675) & comp_A2_124 & comp_A92_250;

assign and_290 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & ~(comp_A92_995) & comp_A996_340 & comp_A998_414;

assign and_291 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & ~(comp_A92_995) & ~(comp_A996_340) & ~(comp_A994_640) & comp_A999_714;

assign and_292 = comp_A93_537 & ~(comp_A9991_972) & ~(comp_A99998_189) & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A99999_594 & ~(comp_A96_754);

assign and_293 = ~(comp_A9991_972) & ~(comp_A9_784) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & comp_A996_332 & comp_A4_484 & comp_A98_325;

assign and_294 = ~(comp_A93_537) & ~(comp_A9991_972) & ~(comp_A92_503) & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & comp_A997_421 & ~(comp_A9996_570);

assign and_295 = ~(comp_A9991_972) & comp_A3_233 & comp_A9_805 & comp_A8_540 & comp_A99996_575;

assign and_296 = ~(comp_A9991_972) & comp_A3_233 & comp_A9_805 & comp_A8_540 & ~(comp_A993_982);

assign and_297 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & ~(comp_A996_332) & comp_A993_659 & ~(comp_A2_602);

assign and_298 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & ~(comp_A996_332) & comp_A993_659 & ~(comp_A92_505);

assign and_299 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & ~(comp_A996_332) & comp_A993_659 & comp_A99999_58;

assign and_300 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & ~(comp_A996_332) & ~(comp_A993_659) & ~(comp_A9992_123);

assign and_301 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A999992_527 & comp_A9996_758 & ~(comp_A997_428) & ~(comp_A93_513) & comp_A99999_558;

assign or_8 = and_274 | and_275 | and_276 | and_277 | and_278 | and_279 | and_280 | and_281 | and_282 | and_283 | and_284 | and_285 | and_286 | and_287 | and_288 | and_289 | and_290 | and_291 | and_292 | and_293 | and_294 | and_295 | and_296 | and_297 | and_298 | and_299 | and_300 | and_301;

assign and_302 = comp_A2_29 & comp_A92_263 & comp_A9991_972 & comp_A1_652 & ~(comp_A991_268) & comp_A99991_539;

assign and_303 = comp_A2_29 & ~(comp_A92_263) & comp_A9991_972 & comp_A1_652 & comp_A7_591;

assign and_304 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & comp_A97_124 & comp_A996_225 & comp_A97_121;

assign and_305 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & ~(comp_A97_124) & comp_A99995_671 & comp_A9998_723;

assign and_306 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & ~(comp_A97_124) & comp_A99995_671 & comp_A999993_9;

assign and_307 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & comp_A997_589 & ~(comp_A97_124) & ~(comp_A99995_671) & ~(comp_A996_92);

assign and_308 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & ~(comp_A996_222) & comp_A91_963;

assign and_309 = ~(comp_A2_29) & comp_A9991_972 & comp_A1_652 & ~(comp_A997_589) & ~(comp_A996_222) & comp_A9994_288;

assign and_310 = ~(comp_A92_263) & comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & ~(comp_A2_901) & comp_A6_406 & comp_A9999_819;

assign and_311 = comp_A9991_972 & ~(comp_A9993_525) & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & ~(comp_A9996_562) & comp_A92_972 & comp_A999995_1015;

assign and_312 = comp_A9991_972 & ~(comp_A995_114) & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & ~(comp_A999996_390) & comp_A92_995 & comp_A996_353 & comp_A99994_600;

assign and_313 = comp_A997_360 & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & comp_A4_486 & comp_A3_232;

assign and_314 = comp_A997_360 & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & ~(comp_A4_486) & comp_A9995_839 & comp_A7_592;

assign and_315 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & comp_A3_286 & comp_A99999_486 & comp_A9991_932;

assign and_316 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & comp_A3_286 & ~(comp_A99999_486) & ~(comp_A996_372);

assign and_317 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & ~(comp_A3_286) & comp_A9_156 & comp_A7_804;

assign and_318 = ~(comp_A997_360) & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & comp_A98_151 & ~(comp_A3_286) & ~(comp_A9_156) & comp_A6_255;

assign and_319 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & comp_A99991_344 & comp_A8_757 & ~(comp_A993_555) & ~(comp_A999994_442);

assign and_320 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & comp_A99991_344 & ~(comp_A8_757) & ~(comp_A99992_671);

assign and_321 = comp_A9992_93 & comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & comp_A99997_931 & ~(comp_A98_151) & ~(comp_A99991_344) & comp_A97_610 & comp_A999991_570;

assign and_322 = comp_A9991_972 & ~(comp_A1_652) & comp_A9991_935 & ~(comp_A99997_931) & ~(comp_A998_424) & comp_A9996_562 & ~(comp_A996_271) & comp_A3_54;

assign and_323 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & comp_A2_901 & comp_A992_675 & ~(comp_A9_821) & comp_A8_536;

assign and_324 = comp_A9991_972 & ~(comp_A1_652) & ~(comp_A9991_935) & ~(comp_A993_317) & comp_A999996_390 & ~(comp_A2_901) & ~(comp_A6_406) & ~(comp_A3_535);

assign and_325 = comp_A93_537 & ~(comp_A9991_972) & comp_A99998_189 & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A99999_594 & ~(comp_A993_492);

assign and_326 = comp_A93_537 & ~(comp_A9991_972) & ~(comp_A99998_189) & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A99999_594 & comp_A96_754;

assign and_327 = ~(comp_A9991_972) & comp_A999992_426 & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & ~(comp_A9996_758) & comp_A9992_429 & ~(comp_A993_440);

assign and_328 = ~(comp_A9991_972) & ~(comp_A9_784) & ~(comp_A3_233) & comp_A9993_530 & comp_A994_475 & comp_A996_332 & ~(comp_A4_484);

assign and_329 = ~(comp_A93_537) & ~(comp_A9991_972) & ~(comp_A3_233) & ~(comp_A9993_530) & comp_A999_712 & ~(comp_A997_421) & ~(comp_A4_445);

assign and_330 = ~(comp_A93_537) & ~(comp_A9991_972) & ~(comp_A3_233) & ~(comp_A9993_530) & ~(comp_A999_712) & comp_A99995_511;

assign and_331 = ~(comp_A9991_972) & comp_A3_233 & ~(comp_A9_805);

assign and_332 = ~(comp_A9991_972) & comp_A3_233 & ~(comp_A8_540);

assign and_333 = ~(comp_A9991_972) & comp_A3_233 & ~(comp_A99996_575) & comp_A993_982;

assign and_334 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & ~(comp_A999992_527);

assign and_335 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & comp_A9996_758 & ~(comp_A997_428) & comp_A93_513;

assign and_336 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & ~(comp_A9996_758) & comp_A9992_429 & comp_A993_440 & comp_A99996_766;

assign and_337 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & ~(comp_A9996_758) & ~(comp_A9992_429) & comp_A999991_485;

assign and_338 = ~(comp_A9991_972) & ~(comp_A3_233) & comp_A9993_530 & ~(comp_A994_475) & ~(comp_A9996_758) & ~(comp_A9992_429) & ~(comp_A9991_1009);

assign or_9 = and_302 | and_303 | and_304 | and_305 | and_306 | and_307 | and_308 | and_309 | and_310 | and_311 | and_312 | and_313 | and_314 | and_315 | and_316 | and_317 | and_318 | and_319 | and_320 | and_321 | and_322 | and_323 | and_324 | and_325 | and_326 | and_327 | and_328 | and_329 | and_330 | and_331 | and_332 | and_333 | and_334 | and_335 | and_336 | and_337 | and_338;

assign and_339 = comp_A3_79 & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & comp_A9991_817;

assign and_340 = comp_A9_827 & ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & ~(comp_A93_651) & ~(comp_A9992_107) & comp_A2_869;

assign and_341 = ~(comp_A4_495) & ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & comp_A3_285 & comp_A94_42 & ~(comp_A97_400);

assign and_342 = comp_A999996_390 & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & ~(comp_A3_305) & comp_A99993_647 & comp_A992_308;

assign and_343 = comp_A99991_185 & comp_A99999_517 & comp_A8_334;

assign and_344 = comp_A99991_185 & comp_A99999_517 & comp_A9996_737 & comp_A9_845 & comp_A997_339 & comp_A997_243 & comp_A993_683;

assign and_345 = comp_A99991_185 & comp_A99999_517 & comp_A9996_737 & comp_A9_845 & comp_A997_339 & ~(comp_A997_243) & ~(comp_A994_543);

assign and_346 = comp_A99991_185 & comp_A99999_517 & ~(comp_A9996_737) & comp_A95_430 & ~(comp_A8_398) & comp_A97_174 & comp_A997_549 & comp_A999996_427;

assign and_347 = comp_A99991_185 & comp_A99999_517 & ~(comp_A9996_737) & comp_A95_430 & ~(comp_A8_398) & ~(comp_A97_174) & comp_A3_381 & comp_A997_496;

assign and_348 = comp_A99991_185 & comp_A99999_517 & ~(comp_A9996_737) & ~(comp_A95_430) & ~(comp_A99_15) & comp_A99_18 & ~(comp_A992_721);

assign and_349 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & comp_A9_853 & ~(comp_A93_136) & ~(comp_A2_320) & comp_A91_383;

assign and_350 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & comp_A9_853 & ~(comp_A93_136) & ~(comp_A2_320) & ~(comp_A6_485);

assign and_351 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & ~(comp_A93_516) & comp_A2_920 & comp_A9991_961 & ~(comp_A999996_360);

assign and_352 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & ~(comp_A93_516) & comp_A2_920 & ~(comp_A9991_961) & ~(comp_A996_350);

assign and_353 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & comp_A96_171 & ~(comp_A98_61);

assign and_354 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & comp_A99996_862 & comp_A9993_327 & ~(comp_A995_537);

assign and_355 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & ~(comp_A99996_862) & ~(comp_A6_442) & comp_A94_58;

assign and_356 = ~(comp_A99991_185) & comp_A99_15 & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & comp_A998_499 & ~(comp_A1_554);

assign and_357 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & comp_A999_567 & ~(comp_A99996_858);

assign and_358 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & comp_A999_567 & comp_A5_316;

assign and_359 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & comp_A999_567 & comp_A995_299;

assign and_360 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & comp_A999_567 & comp_A991_852;

assign and_361 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & ~(comp_A999_567) & comp_A94_49 & comp_A9992_105 & comp_A92_247;

assign and_362 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & ~(comp_A999_567) & comp_A94_49 & ~(comp_A9992_105) & ~(comp_A98_68);

assign and_363 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & ~(comp_A999_567) & ~(comp_A94_49) & ~(comp_A99995_519);

assign and_364 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & comp_A3_285 & comp_A94_42 & comp_A97_400 & ~(comp_A9_155);

assign and_365 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & comp_A3_285 & ~(comp_A94_42) & ~(comp_A3_209);

assign and_366 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & comp_A8_381 & comp_A99_19 & comp_A999997_1011;

assign and_367 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & comp_A998_499 & ~(comp_A1_554) & comp_A999994_662;

assign and_368 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & ~(comp_A998_499) & comp_A5_562 & ~(comp_A9997_669);

assign and_369 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & comp_A9999_248 & comp_A996_245 & ~(comp_A98_1019);

assign and_370 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & comp_A9999_248 & ~(comp_A996_245) & comp_A3_112 & comp_A994_355;

assign and_371 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & comp_A93_651 & comp_A999991_306 & comp_A991_720;

assign and_372 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & ~(comp_A997_578) & comp_A99991_660 & comp_A6_644 & comp_A2_285;

assign and_373 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & ~(comp_A997_578) & ~(comp_A99991_660) & ~(comp_A8_818);

assign and_374 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & comp_A5_505 & comp_A94_35 & comp_A999994_547;

assign and_375 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & comp_A9991_990 & comp_A3_283;

assign or_10 = and_339 | and_340 | and_341 | and_342 | and_343 | and_344 | and_345 | and_346 | and_347 | and_348 | and_349 | and_350 | and_351 | and_352 | and_353 | and_354 | and_355 | and_356 | and_357 | and_358 | and_359 | and_360 | and_361 | and_362 | and_363 | and_364 | and_365 | and_366 | and_367 | and_368 | and_369 | and_370 | and_371 | and_372 | and_373 | and_374 | and_375;

assign and_376 = comp_A9_859 & ~(comp_A999996_390) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & ~(comp_A3_305) & comp_A99993_647;

assign and_377 = ~(comp_A3_79) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & comp_A8_810 & ~(comp_A99994_682) & comp_A9992_99;

assign and_378 = ~(comp_A3_79) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & ~(comp_A8_810) & comp_A9996_610;

assign and_379 = ~(comp_A3_79) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & ~(comp_A8_810) & comp_A997_620;

assign and_380 = comp_A999996_390 & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & ~(comp_A3_305) & comp_A99993_647 & ~(comp_A992_308);

assign and_381 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & comp_A997_339 & ~(comp_A997_243) & comp_A994_543 & comp_A99_13;

assign and_382 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & comp_A2_22 & comp_A92_262 & ~(comp_A96_818);

assign and_383 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & comp_A8_398 & comp_A994_484 & ~(comp_A999997_1009);

assign and_384 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & comp_A8_398 & ~(comp_A994_484) & ~(comp_A3_415);

assign and_385 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & ~(comp_A8_398) & ~(comp_A97_174) & ~(comp_A3_381) & ~(comp_A995_61);

assign and_386 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & ~(comp_A95_430) & comp_A99_15;

assign and_387 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & ~(comp_A95_430) & comp_A99_18 & comp_A992_721 & ~(comp_A6_474);

assign and_388 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & comp_A9_853 & ~(comp_A93_136) & comp_A2_320 & ~(comp_A97_182);

assign and_389 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & comp_A9_853 & ~(comp_A93_136) & ~(comp_A2_320) & ~(comp_A91_383) & comp_A6_485;

assign and_390 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & comp_A93_516 & comp_A99992_501;

assign and_391 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & ~(comp_A93_516) & comp_A2_920 & ~(comp_A9991_961) & comp_A996_350;

assign and_392 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & ~(comp_A93_516) & ~(comp_A2_920) & comp_A991_868 & ~(comp_A992_266);

assign and_393 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & comp_A96_171 & comp_A98_61;

assign and_394 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & comp_A994_378 & comp_A99991_182 & comp_A8_718;

assign and_395 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & comp_A994_378 & ~(comp_A99991_182) & comp_A3_428;

assign and_396 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & comp_A99996_862 & ~(comp_A9993_327) & comp_A9_832;

assign and_397 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & ~(comp_A99996_862) & comp_A6_442 & ~(comp_A999996_428);

assign and_398 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & ~(comp_A99996_862) & ~(comp_A6_442) & ~(comp_A94_58);

assign and_399 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & ~(comp_A9994_693) & comp_A997_521 & comp_A996_360 & comp_A99992_503;

assign and_400 = ~(comp_A99991_185) & ~(comp_A99_15) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & comp_A998_499 & ~(comp_A1_554) & ~(comp_A999994_662);

assign and_401 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & comp_A999_567 & comp_A99996_858 & ~(comp_A5_316) & ~(comp_A995_299) & ~(comp_A991_852);

assign and_402 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & ~(comp_A999_567) & comp_A94_49 & comp_A9992_105 & ~(comp_A92_247);

assign and_403 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & ~(comp_A999_567) & comp_A94_49 & ~(comp_A9992_105) & comp_A98_68;

assign and_404 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & comp_A993_286 & ~(comp_A999_567) & ~(comp_A94_49) & comp_A99995_519;

assign and_405 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & comp_A8_381 & comp_A99_19 & ~(comp_A999997_1011);

assign and_406 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & comp_A8_381 & ~(comp_A99_19) & ~(comp_A92_815);

assign and_407 = comp_A92_264 & ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & ~(comp_A8_381) & comp_A94_33;

assign and_408 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & ~(comp_A998_499) & ~(comp_A5_562);

assign and_409 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & ~(comp_A998_499) & comp_A9997_669 & comp_A997_477;

assign and_410 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & comp_A9999_248 & ~(comp_A996_245) & comp_A3_112 & ~(comp_A994_355) & ~(comp_A993_548);

assign and_411 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & ~(comp_A9999_293) & comp_A92_562 & comp_A99997_252;

assign and_412 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & ~(comp_A9999_293) & comp_A92_562 & comp_A9996_694;

assign and_413 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & comp_A93_651 & ~(comp_A999991_306);

assign and_414 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & comp_A93_651 & ~(comp_A991_720);

assign and_415 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & ~(comp_A93_651) & comp_A9992_107 & comp_A9_851;

assign and_416 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & comp_A997_578 & comp_A998_302;

assign and_417 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & ~(comp_A997_578) & comp_A99991_660 & comp_A6_644 & ~(comp_A2_285);

assign and_418 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & comp_A997_956 & ~(comp_A999992_388) & comp_A991_250 & ~(comp_A95_354);

assign and_419 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & ~(comp_A997_956) & comp_A9994_711 & ~(comp_A9994_295);

assign and_420 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & ~(comp_A5_505) & ~(comp_A9991_956);

assign and_421 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & comp_A9991_990 & ~(comp_A3_283) & comp_A998_641 & ~(comp_A92_377);

assign and_422 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & comp_A9991_990 & ~(comp_A3_283) & ~(comp_A998_641) & ~(comp_A99994_383);

assign and_423 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & comp_A9991_990 & ~(comp_A3_283) & ~(comp_A998_641) & comp_A999992_484;

assign and_424 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & ~(comp_A9991_990) & ~(comp_A9_160) & comp_A997_422;

assign or_11 = and_376 | and_377 | and_378 | and_379 | and_380 | and_381 | and_382 | and_383 | and_384 | and_385 | and_386 | and_387 | and_388 | and_389 | and_390 | and_391 | and_392 | and_393 | and_394 | and_395 | and_396 | and_397 | and_398 | and_399 | and_400 | and_401 | and_402 | and_403 | and_404 | and_405 | and_406 | and_407 | and_408 | and_409 | and_410 | and_411 | and_412 | and_413 | and_414 | and_415 | and_416 | and_417 | and_418 | and_419 | and_420 | and_421 | and_422 | and_423 | and_424;

assign and_425 = ~(comp_A3_79) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & comp_A8_810 & comp_A99994_682 & comp_A993_612;

assign and_426 = ~(comp_A3_79) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & comp_A8_810 & ~(comp_A99994_682) & ~(comp_A9992_99);

assign and_427 = comp_A9_827 & ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & ~(comp_A93_651) & ~(comp_A9992_107) & ~(comp_A2_869);

assign and_428 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & comp_A997_339 & ~(comp_A997_243) & comp_A994_543 & ~(comp_A99_13);

assign and_429 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & ~(comp_A2_22) & comp_A992_528 & ~(comp_A96_271);

assign and_430 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & ~(comp_A2_22) & ~(comp_A992_528) & comp_A994_365;

assign and_431 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & comp_A9_853 & comp_A93_136 & ~(comp_A991_746);

assign and_432 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & ~(comp_A93_516) & comp_A2_920 & comp_A9991_961 & comp_A999996_360;

assign and_433 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & ~(comp_A93_516) & ~(comp_A2_920) & comp_A991_868 & comp_A992_266;

assign and_434 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A99995_471) & ~(comp_A93_516) & ~(comp_A2_920) & ~(comp_A991_868) & ~(comp_A95_312);

assign and_435 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & comp_A994_378 & comp_A99991_182 & ~(comp_A8_718);

assign and_436 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & comp_A994_378 & ~(comp_A99991_182) & ~(comp_A3_428);

assign and_437 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & comp_A99996_862 & comp_A9993_327 & comp_A995_537;

assign and_438 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & ~(comp_A99996_862) & comp_A6_442 & comp_A999996_428;

assign and_439 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & ~(comp_A9994_693) & comp_A997_521 & comp_A996_360 & ~(comp_A99992_503);

assign and_440 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & ~(comp_A8_381) & ~(comp_A94_33) & comp_A9991_937;

assign and_441 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & comp_A997_956 & comp_A999992_388 & ~(comp_A93_687) & ~(comp_A996_292);

assign and_442 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & comp_A5_505 & comp_A94_35 & ~(comp_A999994_547);

assign and_443 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & comp_A5_505 & ~(comp_A94_35) & comp_A9993_685 & comp_A93_718;

assign and_444 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & ~(comp_A5_505) & comp_A9991_956 & comp_A993_484;

assign or_12 = and_425 | and_426 | and_427 | and_428 | and_429 | and_430 | and_431 | and_432 | and_433 | and_434 | and_435 | and_436 | and_437 | and_438 | and_439 | and_440 | and_441 | and_442 | and_443 | and_444;

assign and_445 = comp_A3_79 & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & ~(comp_A9991_817) & comp_A92_246 & comp_A3_27;

assign and_446 = ~(comp_A3_79) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & comp_A8_810 & comp_A99994_682 & ~(comp_A993_612);

assign and_447 = ~(comp_A3_79) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & ~(comp_A8_810) & ~(comp_A9996_610) & ~(comp_A997_620);

assign and_448 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & comp_A2_22 & ~(comp_A92_262) & comp_A3_350;

assign and_449 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & ~(comp_A2_22) & comp_A992_528 & comp_A96_271;

assign and_450 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & ~(comp_A9_845) & comp_A999991_372 & ~(comp_A99999_168);

assign and_451 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & comp_A8_398 & comp_A994_484 & comp_A999997_1009;

assign and_452 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & ~(comp_A8_398) & comp_A97_174 & comp_A997_549 & ~(comp_A999996_427);

assign and_453 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & ~(comp_A8_398) & ~(comp_A97_174) & ~(comp_A3_381) & comp_A995_61;

assign and_454 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & ~(comp_A95_430) & ~(comp_A99_15) & comp_A99_18 & comp_A992_721 & comp_A6_474;

assign and_455 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & comp_A9_853 & comp_A93_136 & comp_A991_746;

assign and_456 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & ~(comp_A9994_693) & comp_A997_521 & ~(comp_A996_360) & ~(comp_A999994_457);

assign and_457 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & ~(comp_A8_381) & ~(comp_A94_33) & ~(comp_A9991_937);

assign and_458 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & comp_A9999_293 & comp_A8_404 & ~(comp_A996_318) & comp_A95_274;

assign and_459 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & comp_A9999_293 & ~(comp_A8_404) & ~(comp_A1_601);

assign and_460 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & ~(comp_A9999_293) & comp_A92_562 & ~(comp_A99997_252) & ~(comp_A9996_694);

assign and_461 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & comp_A3_305 & comp_A997_334 & ~(comp_A999994_507);

assign and_462 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & ~(comp_A997_578) & comp_A99991_660 & ~(comp_A6_644) & comp_A995_202;

assign and_463 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & comp_A997_956 & comp_A999992_388 & comp_A93_687 & comp_A999995_1008;

assign and_464 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & comp_A997_956 & comp_A999992_388 & ~(comp_A93_687) & comp_A996_292;

assign and_465 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & ~(comp_A997_956) & ~(comp_A9994_711);

assign and_466 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & comp_A5_505 & ~(comp_A94_35) & comp_A9993_685 & ~(comp_A93_718);

assign and_467 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & ~(comp_A5_505) & comp_A9991_956 & ~(comp_A993_484) & ~(comp_A1_708);

assign or_13 = and_445 | and_446 | and_447 | and_448 | and_449 | and_450 | and_451 | and_452 | and_453 | and_454 | and_455 | and_456 | and_457 | and_458 | and_459 | and_460 | and_461 | and_462 | and_463 | and_464 | and_465 | and_466 | and_467;

assign and_468 = ~(comp_A9_859) & ~(comp_A999996_390) & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & ~(comp_A3_305);

assign and_469 = comp_A3_79 & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & ~(comp_A9991_817) & ~(comp_A92_246);

assign and_470 = comp_A3_79 & ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & ~(comp_A9999_248) & ~(comp_A9991_817) & ~(comp_A3_27);

assign and_471 = ~(comp_A9_827) & ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & ~(comp_A93_651) & ~(comp_A9992_107);

assign and_472 = comp_A4_495 & ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & comp_A3_285 & comp_A94_42 & ~(comp_A97_400);

assign and_473 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & comp_A997_339 & comp_A997_243 & ~(comp_A993_683);

assign and_474 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & comp_A2_22 & comp_A92_262 & comp_A96_818;

assign and_475 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & comp_A2_22 & ~(comp_A92_262) & ~(comp_A3_350);

assign and_476 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & comp_A9_845 & ~(comp_A997_339) & ~(comp_A2_22) & ~(comp_A992_528) & ~(comp_A994_365);

assign and_477 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & ~(comp_A9_845) & ~(comp_A999991_372);

assign and_478 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & comp_A9996_737 & ~(comp_A9_845) & comp_A99999_168;

assign and_479 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & comp_A8_398 & ~(comp_A994_484) & comp_A3_415;

assign and_480 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & ~(comp_A8_398) & comp_A97_174 & ~(comp_A997_549);

assign and_481 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & comp_A95_430 & ~(comp_A8_398) & ~(comp_A97_174) & comp_A3_381 & ~(comp_A997_496);

assign and_482 = comp_A99991_185 & comp_A99999_517 & ~(comp_A8_334) & ~(comp_A9996_737) & ~(comp_A95_430) & ~(comp_A99_15) & ~(comp_A99_18);

assign and_483 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & ~(comp_A9_853);

assign and_484 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & comp_A2_860 & ~(comp_A93_136) & comp_A2_320 & comp_A97_182;

assign and_485 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & comp_A99995_471;

assign and_486 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & comp_A93_516 & ~(comp_A99992_501);

assign and_487 = comp_A99991_185 & ~(comp_A99999_517) & comp_A95_345 & ~(comp_A2_860) & ~(comp_A93_516) & ~(comp_A2_920) & ~(comp_A991_868) & comp_A95_312;

assign and_488 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & comp_A9994_693 & ~(comp_A994_378) & comp_A99996_862 & ~(comp_A9993_327) & ~(comp_A9_832);

assign and_489 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & ~(comp_A9994_693) & ~(comp_A997_521);

assign and_490 = comp_A99991_185 & ~(comp_A99999_517) & ~(comp_A95_345) & ~(comp_A96_171) & ~(comp_A9994_693) & ~(comp_A996_360) & comp_A999994_457;

assign and_491 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & comp_A3_285 & comp_A94_42 & comp_A97_400 & comp_A9_155;

assign and_492 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & comp_A3_285 & ~(comp_A94_42) & comp_A3_209;

assign and_493 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & comp_A8_381 & ~(comp_A99_19) & comp_A92_815;

assign and_494 = ~(comp_A92_264) & ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & comp_A92_989 & ~(comp_A3_285) & ~(comp_A8_381) & comp_A94_33;

assign and_495 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & comp_A998_499 & comp_A1_554;

assign and_496 = ~(comp_A99991_185) & comp_A99992_710 & comp_A99991_366 & ~(comp_A993_286) & ~(comp_A92_989) & ~(comp_A998_499) & comp_A5_562 & comp_A9997_669 & ~(comp_A997_477);

assign and_497 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & comp_A9999_248 & comp_A996_245 & comp_A98_1019;

assign and_498 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & comp_A9999_248 & ~(comp_A996_245) & ~(comp_A3_112);

assign and_499 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & comp_A9991_973 & comp_A9999_248 & ~(comp_A996_245) & ~(comp_A994_355) & comp_A993_548;

assign and_500 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & comp_A9999_293 & comp_A8_404 & comp_A996_318;

assign and_501 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & comp_A9999_293 & comp_A8_404 & ~(comp_A95_274);

assign and_502 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & comp_A9999_293 & ~(comp_A8_404) & comp_A1_601;

assign and_503 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & comp_A994_477 & ~(comp_A9999_293) & ~(comp_A92_562);

assign and_504 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & comp_A3_305 & ~(comp_A997_334);

assign and_505 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & comp_A3_305 & comp_A999994_507;

assign and_506 = ~(comp_A99991_185) & comp_A99992_710 & ~(comp_A99991_366) & ~(comp_A9991_973) & ~(comp_A994_477) & ~(comp_A3_305) & ~(comp_A99993_647);

assign and_507 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & comp_A997_403 & ~(comp_A93_651) & comp_A9992_107 & ~(comp_A9_851);

assign and_508 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & comp_A997_578 & ~(comp_A998_302);

assign and_509 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & ~(comp_A997_578) & comp_A99991_660 & ~(comp_A6_644) & ~(comp_A995_202);

assign and_510 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & comp_A9993_652 & ~(comp_A997_403) & ~(comp_A997_578) & ~(comp_A99991_660) & comp_A8_818;

assign and_511 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & comp_A997_956 & comp_A999992_388 & comp_A93_687 & ~(comp_A999995_1008);

assign and_512 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & comp_A997_956 & ~(comp_A999992_388) & ~(comp_A991_250);

assign and_513 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & comp_A997_956 & ~(comp_A999992_388) & comp_A95_354;

assign and_514 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & comp_A999995_1012 & ~(comp_A997_956) & comp_A9994_711 & comp_A9994_295;

assign and_515 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & comp_A5_505 & ~(comp_A94_35) & ~(comp_A9993_685);

assign and_516 = ~(comp_A99991_185) & ~(comp_A99992_710) & comp_A99992_810 & ~(comp_A9993_652) & ~(comp_A999995_1012) & ~(comp_A5_505) & comp_A9991_956 & ~(comp_A993_484) & comp_A1_708;

assign and_517 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & comp_A9991_990 & ~(comp_A3_283) & comp_A998_641 & comp_A92_377;

assign and_518 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & comp_A9991_990 & ~(comp_A3_283) & ~(comp_A998_641) & comp_A99994_383 & ~(comp_A999992_484);

assign and_519 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & ~(comp_A9991_990) & comp_A9_160;

assign and_520 = ~(comp_A99991_185) & ~(comp_A99992_710) & ~(comp_A99992_810) & ~(comp_A9991_990) & ~(comp_A997_422);

assign or_14 = and_468 | and_469 | and_470 | and_471 | and_472 | and_473 | and_474 | and_475 | and_476 | and_477 | and_478 | and_479 | and_480 | and_481 | and_482 | and_483 | and_484 | and_485 | and_486 | and_487 | and_488 | and_489 | and_490 | and_491 | and_492 | and_493 | and_494 | and_495 | and_496 | and_497 | and_498 | and_499 | and_500 | and_501 | and_502 | and_503 | and_504 | and_505 | and_506 | and_507 | and_508 | and_509 | and_510 | and_511 | and_512 | and_513 | and_514 | and_515 | and_516 | and_517 | and_518 | and_519 | and_520;

assign and_521 = comp_A98_171 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & ~(comp_A9996_693) & ~(comp_A99996_513);

assign and_522 = ~(comp_A94_46) & comp_A9_827 & comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A2_827 & comp_A999997_1012;

assign and_523 = comp_A999997_1009 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & comp_A999_585 & ~(comp_A5_753) & comp_A7_856;

assign and_524 = comp_A99991_182 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & comp_A997_666 & ~(comp_A94_37) & comp_A996_343;

assign and_525 = comp_A2_862 & comp_A96_180 & comp_A99997_843 & comp_A9994_704 & comp_A98_240;

assign and_526 = comp_A2_862 & comp_A96_180 & comp_A99997_843 & ~(comp_A9994_704) & ~(comp_A3_992);

assign and_527 = comp_A94_46 & comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A2_827 & comp_A999997_1012 & comp_A994_549;

assign and_528 = comp_A94_46 & comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A2_827 & comp_A999997_1012 & ~(comp_A97_171);

assign and_529 = ~(comp_A94_46) & comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A2_827 & comp_A999997_1012 & comp_A9993_313;

assign and_530 = comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A2_827 & ~(comp_A999997_1012) & ~(comp_A4_545);

assign and_531 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & comp_A93_115 & comp_A9991_962 & comp_A99993_596;

assign and_532 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & comp_A2_114 & comp_A995_493 & comp_A99996_188 & comp_A3_116;

assign and_533 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & comp_A2_114 & ~(comp_A995_493) & ~(comp_A2_9);

assign and_534 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & comp_A2_114 & ~(comp_A995_493) & comp_A93_544;

assign and_535 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & ~(comp_A2_114) & comp_A3_812 & comp_A997_373;

assign and_536 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & ~(comp_A2_114) & ~(comp_A3_812) & comp_A9991_955 & comp_A9998_906;

assign and_537 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & comp_A999_585 & comp_A5_753 & ~(comp_A99993_51) & ~(comp_A92_255);

assign and_538 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & ~(comp_A999_585) & comp_A9_829 & comp_A99995_559 & ~(comp_A2_33);

assign and_539 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & ~(comp_A997_666) & comp_A996_263 & ~(comp_A9996_763) & ~(comp_A99992_660);

assign and_540 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & comp_A997_381 & comp_A99992_538;

assign and_541 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & ~(comp_A97_201) & comp_A994_677 & comp_A99_18 & ~(comp_A93_720);

assign and_542 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & comp_A996_244 & ~(comp_A9999_786) & comp_A97_968 & comp_A9993_626;

assign and_543 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & comp_A996_244 & ~(comp_A9999_786) & ~(comp_A97_968) & comp_A99998_187;

assign and_544 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & comp_A92_528 & ~(comp_A7_460) & ~(comp_A98_153) & ~(comp_A999_516);

assign and_545 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & comp_A991_373 & comp_A9993_658 & ~(comp_A999992_474) & comp_A999995_1014;

assign or_15 = and_521 | and_522 | and_523 | and_524 | and_525 | and_526 | and_527 | and_528 | and_529 | and_530 | and_531 | and_532 | and_533 | and_534 | and_535 | and_536 | and_537 | and_538 | and_539 | and_540 | and_541 | and_542 | and_543 | and_544 | and_545;

assign and_546 = ~(comp_A98_171) & comp_A92_503 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & comp_A997_451;

assign and_547 = ~(comp_A94_46) & ~(comp_A9_827) & comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A999997_1012 & ~(comp_A9993_313);

assign and_548 = ~(comp_A9_156) & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & comp_A92_528 & comp_A7_460 & ~(comp_A93_722);

assign and_549 = comp_A2_920 & ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & comp_A97_201 & ~(comp_A3_750);

assign and_550 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & comp_A996_327 & comp_A1_684 & comp_A99999_443;

assign and_551 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & comp_A996_327 & ~(comp_A1_684) & comp_A9996_623;

assign and_552 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & ~(comp_A996_327) & ~(comp_A9_150) & ~(comp_A9991_965);

assign and_553 = ~(comp_A99992_810) & ~(comp_A999995_1008) & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & ~(comp_A999992_432);

assign and_554 = ~(comp_A99992_810) & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & ~(comp_A999992_432) & ~(comp_A999996_726);

assign and_555 = comp_A9992_103 & ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & comp_A997_381 & ~(comp_A99992_538) & ~(comp_A99994_755);

assign and_556 = comp_A2_862 & comp_A96_180 & comp_A99997_843 & comp_A9994_704 & ~(comp_A98_240);

assign and_557 = comp_A2_862 & comp_A96_180 & comp_A99997_843 & ~(comp_A9994_704) & comp_A3_992 & comp_A9994_881;

assign and_558 = comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & ~(comp_A2_827);

assign and_559 = comp_A94_46 & comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A999997_1012 & ~(comp_A994_549) & comp_A97_171;

assign and_560 = comp_A2_862 & ~(comp_A96_180) & comp_A996_200 & ~(comp_A3_247) & comp_A995_185 & ~(comp_A998_559) & ~(comp_A9999_767);

assign and_561 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & comp_A93_115 & comp_A9991_962 & ~(comp_A99993_596) & ~(comp_A93_98);

assign and_562 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & comp_A93_115 & ~(comp_A9991_962) & comp_A99994_807 & ~(comp_A96_264);

assign and_563 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & comp_A93_115 & ~(comp_A9991_962) & ~(comp_A99994_807) & comp_A92_500;

assign and_564 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & comp_A2_114 & comp_A995_493 & ~(comp_A99996_188) & comp_A99996_839;

assign and_565 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & comp_A2_114 & ~(comp_A995_493) & comp_A2_9 & ~(comp_A93_544);

assign and_566 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & ~(comp_A2_114) & comp_A3_812 & ~(comp_A997_373) & ~(comp_A99999_423);

assign and_567 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & ~(comp_A2_114) & ~(comp_A3_812) & ~(comp_A9991_955);

assign and_568 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & comp_A997_666 & comp_A94_37 & ~(comp_A9991_1011) & ~(comp_A99991_408);

assign and_569 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & comp_A997_666 & ~(comp_A94_37) & ~(comp_A996_343) & ~(comp_A9999_560);

assign and_570 = ~(comp_A2_862) & comp_A1_642 & ~(comp_A9999_419) & ~(comp_A7_643) & ~(comp_A99992_736);

assign and_571 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & ~(comp_A997_381) & ~(comp_A99992_655) & comp_A3_386 & comp_A9998_389;

assign and_572 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & ~(comp_A997_381) & ~(comp_A99992_655) & ~(comp_A3_386) & ~(comp_A994_390);

assign and_573 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & comp_A97_201 & ~(comp_A3_750) & comp_A995_34;

assign and_574 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & ~(comp_A97_201) & comp_A994_677 & ~(comp_A99_18) & comp_A99997_149;

assign and_575 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & comp_A996_244 & comp_A9999_786 & ~(comp_A99992_744);

assign and_576 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & comp_A996_244 & ~(comp_A9999_786) & comp_A97_968 & ~(comp_A9993_626);

assign and_577 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & comp_A996_244 & ~(comp_A9999_786) & ~(comp_A97_968) & ~(comp_A99998_187);

assign and_578 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & ~(comp_A996_244) & comp_A99994_612 & comp_A9991_982 & comp_A2_918;

assign and_579 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & ~(comp_A996_244) & comp_A99994_612 & ~(comp_A9991_982) & ~(comp_A996_304);

assign and_580 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & ~(comp_A996_244) & ~(comp_A99994_612) & comp_A99_5 & ~(comp_A9991_693);

assign and_581 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & ~(comp_A996_244) & ~(comp_A99994_612) & ~(comp_A99_5) & ~(comp_A99_21);

assign and_582 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & comp_A3_103 & comp_A998_676 & ~(comp_A9_486);

assign and_583 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & comp_A991_373 & comp_A9993_658 & comp_A999992_474;

assign and_584 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & comp_A991_373 & comp_A9993_658 & ~(comp_A999995_1014);

assign and_585 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & comp_A991_373 & ~(comp_A9993_658) & ~(comp_A9995_441);

assign or_16 = and_546 | and_547 | and_548 | and_549 | and_550 | and_551 | and_552 | and_553 | and_554 | and_555 | and_556 | and_557 | and_558 | and_559 | and_560 | and_561 | and_562 | and_563 | and_564 | and_565 | and_566 | and_567 | and_568 | and_569 | and_570 | and_571 | and_572 | and_573 | and_574 | and_575 | and_576 | and_577 | and_578 | and_579 | and_580 | and_581 | and_582 | and_583 | and_584 | and_585;

assign and_586 = comp_A98_171 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & comp_A9996_693 & comp_A99993_630;

assign and_587 = comp_A9_156 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & comp_A92_528 & comp_A7_460 & comp_A999994_411;

assign and_588 = ~(comp_A9_156) & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & comp_A92_528 & comp_A7_460 & comp_A93_722;

assign and_589 = comp_A999997_1009 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & comp_A999_585 & ~(comp_A5_753) & ~(comp_A7_856);

assign and_590 = ~(comp_A2_920) & ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & comp_A97_201 & ~(comp_A3_750) & ~(comp_A995_34);

assign and_591 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & ~(comp_A996_327) & ~(comp_A9_150) & comp_A9991_965;

assign and_592 = ~(comp_A9992_103) & ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & comp_A997_381 & ~(comp_A99992_538) & ~(comp_A99994_755);

assign and_593 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & comp_A93_115 & ~(comp_A9991_962) & ~(comp_A99994_807) & ~(comp_A92_500);

assign and_594 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & ~(comp_A999_585) & comp_A9_829 & comp_A99995_559 & comp_A2_33;

assign and_595 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & ~(comp_A999_585) & ~(comp_A9_829) & comp_A9992_436;

assign and_596 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & ~(comp_A997_666) & comp_A996_263 & ~(comp_A9996_763) & comp_A99992_660;

assign and_597 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & ~(comp_A997_381) & comp_A99992_655 & ~(comp_A991_451) & comp_A99995_531;

assign and_598 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & ~(comp_A997_381) & ~(comp_A99992_655) & ~(comp_A3_386) & comp_A994_390;

assign and_599 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & ~(comp_A996_244) & ~(comp_A99994_612) & comp_A99_5 & comp_A9991_693;

assign and_600 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A9_151) & ~(comp_A996_244) & ~(comp_A99994_612) & ~(comp_A99_5) & comp_A99_21;

assign and_601 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & comp_A92_528 & ~(comp_A7_460) & comp_A98_153 & comp_A996_231;

assign or_17 = and_586 | and_587 | and_588 | and_589 | and_590 | and_591 | and_592 | and_593 | and_594 | and_595 | and_596 | and_597 | and_598 | and_599 | and_600 | and_601;

assign and_602 = comp_A98_171 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & ~(comp_A9996_693) & comp_A99996_513;

assign and_603 = ~(comp_A98_171) & ~(comp_A92_503) & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & comp_A9992_161;

assign and_604 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & ~(comp_A996_327) & comp_A9_150 & ~(comp_A997_713);

assign and_605 = comp_A2_862 & ~(comp_A96_180) & comp_A996_200 & ~(comp_A3_247) & comp_A995_185 & ~(comp_A998_559) & comp_A9999_767;

assign and_606 = comp_A2_862 & ~(comp_A96_180) & comp_A996_200 & ~(comp_A3_247) & ~(comp_A995_185) & ~(comp_A99996_551);

assign and_607 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & comp_A93_115 & comp_A9991_962 & ~(comp_A99993_596) & comp_A93_98;

assign and_608 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & comp_A2_114 & comp_A995_493 & comp_A99996_188 & ~(comp_A3_116);

assign and_609 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & ~(comp_A999_585) & comp_A9_829 & ~(comp_A99995_559) & ~(comp_A99999_545);

assign and_610 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & ~(comp_A997_666) & ~(comp_A996_263);

assign and_611 = ~(comp_A2_862) & comp_A1_642 & ~(comp_A9999_419) & ~(comp_A7_643) & comp_A99992_736 & ~(comp_A9_61);

assign and_612 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & comp_A997_381 & ~(comp_A99992_538) & comp_A99994_755 & ~(comp_A8_484);

assign and_613 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & comp_A97_201 & comp_A3_750;

assign and_614 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & ~(comp_A97_201) & comp_A994_677 & comp_A99_18 & comp_A93_720;

assign and_615 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & ~(comp_A97_201) & ~(comp_A994_677) & comp_A3_588;

assign and_616 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & ~(comp_A97_201) & ~(comp_A994_677) & ~(comp_A98_120);

assign and_617 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & comp_A92_528 & ~(comp_A7_460) & comp_A98_153 & ~(comp_A996_231);

assign or_18 = and_602 | and_603 | and_604 | and_605 | and_606 | and_607 | and_608 | and_609 | and_610 | and_611 | and_612 | and_613 | and_614 | and_615 | and_616 | and_617;

assign and_618 = comp_A98_171 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & comp_A9996_693 & ~(comp_A99993_630);

assign and_619 = ~(comp_A98_171) & comp_A92_503 & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & ~(comp_A997_451);

assign and_620 = ~(comp_A98_171) & ~(comp_A92_503) & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & ~(comp_A93_115) & ~(comp_A9992_161);

assign and_621 = comp_A9_156 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & comp_A7_460 & ~(comp_A999994_411);

assign and_622 = ~(comp_A999997_1009) & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & comp_A999_585 & ~(comp_A5_753);

assign and_623 = ~(comp_A99991_182) & comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & comp_A997_666 & ~(comp_A94_37) & comp_A996_343;

assign and_624 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & comp_A996_327 & comp_A1_684 & ~(comp_A99999_443);

assign and_625 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & comp_A996_327 & ~(comp_A1_684) & ~(comp_A9996_623);

assign and_626 = comp_A99992_810 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & ~(comp_A996_327) & comp_A9_150 & comp_A997_713;

assign and_627 = ~(comp_A99992_810) & comp_A999995_1008 & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & comp_A999996_726;

assign and_628 = ~(comp_A99992_810) & ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & ~(comp_A991_373) & comp_A999992_432;

assign and_629 = comp_A2_862 & comp_A96_180 & comp_A99997_843 & ~(comp_A9994_704) & comp_A3_992 & ~(comp_A9994_881);

assign and_630 = comp_A2_862 & comp_A96_180 & ~(comp_A99997_843) & comp_A2_827 & ~(comp_A999997_1012) & comp_A4_545;

assign and_631 = comp_A2_862 & ~(comp_A96_180) & comp_A996_200 & comp_A3_247;

assign and_632 = comp_A2_862 & ~(comp_A96_180) & comp_A996_200 & comp_A995_185 & comp_A998_559;

assign and_633 = comp_A2_862 & ~(comp_A96_180) & comp_A996_200 & ~(comp_A995_185) & comp_A99996_551;

assign and_634 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & comp_A992_817 & comp_A93_115 & ~(comp_A9991_962) & comp_A99994_807 & comp_A96_264;

assign and_635 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & comp_A2_114 & comp_A995_493 & ~(comp_A99996_188) & ~(comp_A99996_839);

assign and_636 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & ~(comp_A2_114) & comp_A3_812 & ~(comp_A997_373) & comp_A99999_423;

assign and_637 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & comp_A6_701 & ~(comp_A992_817) & ~(comp_A2_114) & ~(comp_A3_812) & comp_A9991_955 & ~(comp_A9998_906);

assign and_638 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & comp_A999_585 & comp_A5_753 & comp_A99993_51;

assign and_639 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & comp_A999_585 & comp_A5_753 & comp_A92_255;

assign and_640 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & ~(comp_A999_585) & comp_A9_829 & ~(comp_A99995_559) & comp_A99999_545;

assign and_641 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & comp_A999996_461 & ~(comp_A999_585) & ~(comp_A9_829) & ~(comp_A9992_436);

assign and_642 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & comp_A997_666 & comp_A94_37 & comp_A9991_1011;

assign and_643 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & comp_A997_666 & comp_A94_37 & comp_A99991_408;

assign and_644 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & comp_A997_666 & ~(comp_A94_37) & ~(comp_A996_343) & comp_A9999_560;

assign and_645 = comp_A2_862 & ~(comp_A96_180) & ~(comp_A996_200) & ~(comp_A6_701) & ~(comp_A999996_461) & ~(comp_A997_666) & comp_A996_263 & comp_A9996_763;

assign and_646 = ~(comp_A2_862) & comp_A1_642 & comp_A9999_419;

assign and_647 = ~(comp_A2_862) & comp_A1_642 & comp_A7_643;

assign and_648 = ~(comp_A2_862) & comp_A1_642 & comp_A99992_736 & comp_A9_61;

assign and_649 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & comp_A997_381 & ~(comp_A99992_538) & comp_A99994_755 & comp_A8_484;

assign and_650 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & ~(comp_A997_381) & comp_A99992_655 & comp_A991_451;

assign and_651 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & ~(comp_A997_381) & comp_A99992_655 & ~(comp_A99995_531);

assign and_652 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & comp_A3_565 & ~(comp_A997_381) & ~(comp_A99992_655) & comp_A3_386 & ~(comp_A9998_389);

assign and_653 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & ~(comp_A97_201) & comp_A994_677 & ~(comp_A99_18) & ~(comp_A99997_149);

assign and_654 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & comp_A99999_406 & ~(comp_A3_565) & ~(comp_A97_201) & ~(comp_A994_677) & ~(comp_A3_588) & comp_A98_120;

assign and_655 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & comp_A9_151;

assign and_656 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & comp_A996_244 & comp_A9999_786 & comp_A99992_744;

assign and_657 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A996_244) & comp_A99994_612 & comp_A9991_982 & ~(comp_A2_918);

assign and_658 = ~(comp_A2_862) & ~(comp_A1_642) & comp_A6_394 & ~(comp_A99999_406) & ~(comp_A996_244) & comp_A99994_612 & ~(comp_A9991_982) & comp_A996_304;

assign and_659 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & comp_A3_103 & ~(comp_A998_676);

assign and_660 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & comp_A3_103 & comp_A9_486;

assign and_661 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & ~(comp_A92_528);

assign and_662 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & comp_A9991_931 & ~(comp_A3_103) & ~(comp_A7_460) & ~(comp_A98_153) & comp_A999_516;

assign and_663 = ~(comp_A2_862) & ~(comp_A1_642) & ~(comp_A6_394) & ~(comp_A9991_931) & comp_A991_373 & ~(comp_A9993_658) & comp_A9995_441;

assign or_19 = and_618 | and_619 | and_620 | and_621 | and_622 | and_623 | and_624 | and_625 | and_626 | and_627 | and_628 | and_629 | and_630 | and_631 | and_632 | and_633 | and_634 | and_635 | and_636 | and_637 | and_638 | and_639 | and_640 | and_641 | and_642 | and_643 | and_644 | and_645 | and_646 | and_647 | and_648 | and_649 | and_650 | and_651 | and_652 | and_653 | and_654 | and_655 | and_656 | and_657 | and_658 | and_659 | and_660 | and_661 | and_662 | and_663;

assign and_664 = ~(comp_A97_193) & comp_A3_79 & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955;

assign and_665 = ~(comp_A97_193) & comp_A9_811 & ~(comp_A92_995) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & ~(comp_A93_92);

assign and_666 = ~(comp_A97_193) & ~(comp_A9_811) & ~(comp_A92_995) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & comp_A9991_932;

assign and_667 = comp_A97_193 & ~(comp_A92_246) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & ~(comp_A999996_685) & comp_A99992_711 & ~(comp_A9991_921);

assign and_668 = comp_A97_193 & ~(comp_A9_150) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & comp_A999996_685 & ~(comp_A2_844) & comp_A991_391;

assign and_669 = comp_A97_193 & comp_A993_258;

assign and_670 = comp_A97_193 & comp_A8_335 & comp_A999_656;

assign and_671 = comp_A97_193 & comp_A8_335 & comp_A991_735;

assign and_672 = comp_A97_193 & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & comp_A999996_685 & comp_A2_844 & comp_A997_399;

assign and_673 = ~(comp_A97_193) & comp_A9_816 & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & comp_A93_119 & comp_A992_234 & comp_A92_992;

assign and_674 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & ~(comp_A1_581) & comp_A993_621 & ~(comp_A999992_339) & ~(comp_A99993_85);

assign and_675 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & comp_A93_119 & comp_A992_234 & ~(comp_A92_992) & ~(comp_A991_644);

assign and_676 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & ~(comp_A996_311) & comp_A997_299 & comp_A99992_670;

assign and_677 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & comp_A1_741 & comp_A994_524 & comp_A9997_340;

assign and_678 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & comp_A1_741 & ~(comp_A994_524) & ~(comp_A99994_727) & comp_A994_644;

assign and_679 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & comp_A3_127 & ~(comp_A6_452) & ~(comp_A4_332);

assign and_680 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & ~(comp_A3_127) & comp_A8_875 & comp_A97_207 & ~(comp_A9993_671);

assign or_20 = and_664 | and_665 | and_666 | and_667 | and_668 | and_669 | and_670 | and_671 | and_672 | and_673 | and_674 | and_675 | and_676 | and_677 | and_678 | and_679 | and_680;

assign and_681 = ~(comp_A97_193) & ~(comp_A3_79) & ~(comp_A9_811) & ~(comp_A92_995) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & ~(comp_A9991_932);

assign and_682 = ~(comp_A97_193) & ~(comp_A3_79) & comp_A92_995 & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & comp_A991_647 & ~(comp_A996_185);

assign and_683 = comp_A97_193 & ~(comp_A92_246) & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & ~(comp_A999996_685) & ~(comp_A99992_711);

assign and_684 = comp_A97_193 & ~(comp_A92_246) & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & ~(comp_A999996_685) & comp_A9991_921;

assign and_685 = comp_A97_193 & ~(comp_A993_258) & comp_A8_335 & ~(comp_A999_656) & ~(comp_A991_735);

assign and_686 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & comp_A996_203 & comp_A93_546 & comp_A99996_508 & ~(comp_A99996_263);

assign and_687 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & comp_A94_30 & comp_A999_711 & comp_A9_840 & ~(comp_A91_210);

assign and_688 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & comp_A94_30 & comp_A999_711 & comp_A9_840 & comp_A9997_587;

assign and_689 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & comp_A94_30 & ~(comp_A999_711) & ~(comp_A2_713);

assign and_690 = ~(comp_A97_193) & ~(comp_A9_816) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & comp_A93_119 & comp_A992_234 & comp_A92_992;

assign and_691 = ~(comp_A97_193) & ~(comp_A9_821) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & comp_A93_119 & ~(comp_A992_234);

assign and_692 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & ~(comp_A1_581) & comp_A993_621 & ~(comp_A999992_339) & comp_A99993_85;

assign and_693 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & comp_A93_119 & comp_A992_234 & ~(comp_A92_992) & comp_A991_644;

assign and_694 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & comp_A93_119 & ~(comp_A992_234) & comp_A3_662;

assign and_695 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & ~(comp_A996_311) & comp_A997_299 & ~(comp_A99992_670);

assign and_696 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & ~(comp_A996_311) & ~(comp_A997_299) & comp_A94_32;

assign and_697 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & comp_A1_741 & ~(comp_A994_524) & ~(comp_A99994_727) & ~(comp_A994_644);

assign and_698 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & comp_A996_369 & comp_A9991_995 & comp_A5_492;

assign and_699 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & comp_A996_369 & ~(comp_A9991_995) & ~(comp_A998_230);

assign and_700 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & ~(comp_A996_369) & ~(comp_A93_532) & comp_A95_388;

assign and_701 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & comp_A3_127 & comp_A6_452;

assign and_702 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & comp_A3_127 & comp_A4_332 & comp_A999996_581;

assign and_703 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & ~(comp_A3_127) & ~(comp_A8_875) & comp_A9991_699;

assign or_21 = and_681 | and_682 | and_683 | and_684 | and_685 | and_686 | and_687 | and_688 | and_689 | and_690 | and_691 | and_692 | and_693 | and_694 | and_695 | and_696 | and_697 | and_698 | and_699 | and_700 | and_701 | and_702 | and_703;

assign and_704 = ~(comp_A97_193) & ~(comp_A3_79) & comp_A92_995 & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & ~(comp_A991_647) & comp_A999992_536;

assign and_705 = comp_A97_193 & ~(comp_A9_150) & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & comp_A999996_685 & ~(comp_A2_844) & ~(comp_A991_391);

assign and_706 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & comp_A94_30 & comp_A999_711 & comp_A9_840 & comp_A91_210 & ~(comp_A9997_587);

assign and_707 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & comp_A999996_685 & comp_A2_844 & ~(comp_A997_399) & comp_A9993_561;

assign and_708 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & comp_A1_581 & ~(comp_A991_486);

assign and_709 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & ~(comp_A1_581) & ~(comp_A993_621) & comp_A92_574 & comp_A3_867;

assign and_710 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & comp_A996_311 & comp_A994_457 & comp_A9993_539;

assign and_711 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & comp_A3_127 & ~(comp_A6_452) & comp_A4_332 & ~(comp_A999996_581);

assign or_22 = and_704 | and_705 | and_706 | and_707 | and_708 | and_709 | and_710 | and_711;

assign and_712 = ~(comp_A97_193) & ~(comp_A3_79) & comp_A9_811 & ~(comp_A92_995) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & comp_A93_92;

assign and_713 = ~(comp_A97_193) & ~(comp_A3_79) & comp_A92_995 & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & comp_A991_647 & comp_A996_185;

assign and_714 = comp_A97_193 & comp_A92_246 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & ~(comp_A999996_685) & ~(comp_A6_286);

assign and_715 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & comp_A996_203 & comp_A93_546 & ~(comp_A99996_508);

assign and_716 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & comp_A996_203 & ~(comp_A93_546) & ~(comp_A9996_431) & comp_A96_22;

assign and_717 = ~(comp_A97_193) & comp_A9_821 & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & comp_A93_119 & ~(comp_A992_234) & ~(comp_A3_662);

assign and_718 = ~(comp_A97_193) & comp_A92_246 & comp_A99995_531 & comp_A3_55 & ~(comp_A9_157) & comp_A991_797 & comp_A997_394 & comp_A96_766 & comp_A9993_581;

assign and_719 = ~(comp_A97_193) & comp_A92_246 & comp_A3_55 & comp_A9_157 & comp_A8_657 & comp_A99994_586;

assign and_720 = ~(comp_A97_193) & comp_A92_246 & comp_A3_55 & ~(comp_A9_157) & ~(comp_A991_797) & comp_A9998_661;

assign and_721 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & comp_A1_581 & comp_A991_486;

assign and_722 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & ~(comp_A1_581) & comp_A993_621 & comp_A999992_339 & ~(comp_A7_767);

assign and_723 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & ~(comp_A1_581) & ~(comp_A993_621) & comp_A92_574 & ~(comp_A3_867);

assign and_724 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & comp_A996_311 & ~(comp_A994_457) & ~(comp_A99997_946);

assign and_725 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & ~(comp_A996_311) & ~(comp_A997_299) & ~(comp_A94_32);

assign and_726 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & comp_A1_741 & comp_A994_524 & ~(comp_A9997_340) & ~(comp_A997_696);

assign and_727 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & ~(comp_A996_369) & comp_A93_532 & comp_A999_337;

assign and_728 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & ~(comp_A3_127) & comp_A8_875 & ~(comp_A97_207) & comp_A9999_59 & ~(comp_A991_777);

assign or_23 = and_712 | and_713 | and_714 | and_715 | and_716 | and_717 | and_718 | and_719 | and_720 | and_721 | and_722 | and_723 | and_724 | and_725 | and_726 | and_727 | and_728;

assign and_729 = ~(comp_A97_193) & ~(comp_A3_79) & comp_A92_995 & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & comp_A99997_955 & ~(comp_A991_647) & ~(comp_A999992_536);

assign and_730 = comp_A97_193 & comp_A92_246 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & ~(comp_A999996_685) & comp_A6_286;

assign and_731 = comp_A97_193 & comp_A9_150 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & comp_A999996_685 & ~(comp_A2_844);

assign and_732 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & comp_A996_203 & comp_A93_546 & comp_A99996_508 & comp_A99996_263;

assign and_733 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & comp_A996_203 & ~(comp_A93_546) & comp_A9996_431;

assign and_734 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & comp_A996_203 & ~(comp_A93_546) & ~(comp_A96_22);

assign and_735 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & comp_A94_30 & comp_A999_711 & ~(comp_A9_840);

assign and_736 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & comp_A94_30 & ~(comp_A999_711) & comp_A2_713;

assign and_737 = comp_A97_193 & ~(comp_A993_258) & ~(comp_A8_335) & ~(comp_A996_203) & ~(comp_A94_30) & comp_A999996_685 & comp_A2_844 & ~(comp_A997_399) & ~(comp_A9993_561);

assign and_738 = ~(comp_A97_193) & ~(comp_A92_246) & comp_A3_55;

assign and_739 = ~(comp_A97_193) & ~(comp_A99995_531) & comp_A3_55 & ~(comp_A9_157) & comp_A991_797;

assign and_740 = ~(comp_A97_193) & comp_A3_55 & comp_A9_157 & ~(comp_A8_657);

assign and_741 = ~(comp_A97_193) & comp_A3_55 & comp_A9_157 & ~(comp_A99994_586);

assign and_742 = ~(comp_A97_193) & comp_A3_55 & ~(comp_A9_157) & comp_A991_797 & ~(comp_A997_394);

assign and_743 = ~(comp_A97_193) & comp_A3_55 & ~(comp_A9_157) & comp_A991_797 & ~(comp_A96_766);

assign and_744 = ~(comp_A97_193) & comp_A3_55 & ~(comp_A9_157) & comp_A991_797 & ~(comp_A9993_581);

assign and_745 = ~(comp_A97_193) & comp_A3_55 & ~(comp_A9_157) & ~(comp_A991_797) & ~(comp_A9998_661);

assign and_746 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & ~(comp_A1_581) & comp_A993_621 & comp_A999992_339 & comp_A7_767;

assign and_747 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & comp_A9996_707 & ~(comp_A99997_955) & ~(comp_A1_581) & ~(comp_A993_621) & ~(comp_A92_574);

assign and_748 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & comp_A996_311 & comp_A994_457 & ~(comp_A9993_539);

assign and_749 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & comp_A98_270 & ~(comp_A93_119) & comp_A996_311 & ~(comp_A994_457) & comp_A99997_946;

assign and_750 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & comp_A1_741 & comp_A994_524 & ~(comp_A9997_340) & comp_A997_696;

assign and_751 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & comp_A1_741 & ~(comp_A994_524) & comp_A99994_727;

assign and_752 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & comp_A996_369 & comp_A9991_995 & ~(comp_A5_492);

assign and_753 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & comp_A996_369 & ~(comp_A9991_995) & comp_A998_230;

assign and_754 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & ~(comp_A996_369) & comp_A93_532 & ~(comp_A999_337);

assign and_755 = ~(comp_A97_193) & ~(comp_A3_55) & comp_A99993_699 & ~(comp_A9996_707) & ~(comp_A98_270) & ~(comp_A1_741) & ~(comp_A996_369) & ~(comp_A93_532) & ~(comp_A95_388);

assign and_756 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & ~(comp_A3_127) & comp_A8_875 & comp_A97_207 & comp_A9993_671;

assign and_757 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & ~(comp_A3_127) & comp_A8_875 & ~(comp_A97_207) & ~(comp_A9999_59);

assign and_758 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & ~(comp_A3_127) & comp_A8_875 & ~(comp_A97_207) & comp_A991_777;

assign and_759 = ~(comp_A97_193) & ~(comp_A3_55) & ~(comp_A99993_699) & ~(comp_A3_127) & ~(comp_A8_875) & ~(comp_A9991_699);

assign or_24 = and_729 | and_730 | and_731 | and_732 | and_733 | and_734 | and_735 | and_736 | and_737 | and_738 | and_739 | and_740 | and_741 | and_742 | and_743 | and_744 | and_745 | and_746 | and_747 | and_748 | and_749 | and_750 | and_751 | and_752 | and_753 | and_754 | and_755 | and_756 | and_757 | and_758 | and_759;


endmodule


module MAJ(
or_0, or_1, or_2, or_3, or_4, or_5, or_6, or_7, or_8, or_9, or_10, or_11, or_12, or_13, or_14, or_15, or_16, or_17, or_18, or_19, or_20, or_21, or_22, or_23, or_24, reg_decision
);

input [0:0] or_0;
input [0:0] or_1;
input [0:0] or_2;
input [0:0] or_3;
input [0:0] or_4;
input [0:0] or_5;
input [0:0] or_6;
input [0:0] or_7;
input [0:0] or_8;
input [0:0] or_9;
input [0:0] or_10;
input [0:0] or_11;
input [0:0] or_12;
input [0:0] or_13;
input [0:0] or_14;
input [0:0] or_15;
input [0:0] or_16;
input [0:0] or_17;
input [0:0] or_18;
input [0:0] or_19;
input [0:0] or_20;
input [0:0] or_21;
input [0:0] or_22;
input [0:0] or_23;
input [0:0] or_24;
output [4:0] reg_decision;
wire [2:0] add_0;
wire [2:0] add_1;
wire [2:0] add_2;
wire [2:0] add_3;
wire [2:0] add_4;
wire [0:0] comp_add_0_1;
wire [0:0] comp_add_2_3;
wire [0:0] comp_add_0_1_2_3;
wire [0:0] comp_add_0_1_2_3_4;
wire [2:0] add_0_1;
wire [2:0] add_2_3;
wire [2:0] add_0_1_2_3;
wire [2:0] add_0_1_2_3_4;
wire [2:0] sel_decision_0;
wire [2:0] sel_decision_1;
wire [2:0] sel_decision_2;
wire [2:0] sel_decision_3;
wire [0:0] sel_decision_4;

assign add_0 = {2'b00, or_0} + {2'b00, or_5} + {2'b00, or_10} + {2'b00, or_15} + {2'b00, or_20};

assign add_1 = {2'b00, or_1} + {2'b00, or_6} + {2'b00, or_11} + {2'b00, or_16} + {2'b00, or_21};

assign add_2 = {2'b00, or_2} + {2'b00, or_7} + {2'b00, or_12} + {2'b00, or_17} + {2'b00, or_22};

assign add_3 = {2'b00, or_3} + {2'b00, or_8} + {2'b00, or_13} + {2'b00, or_18} + {2'b00, or_23};

assign add_4 = {2'b00, or_4} + {2'b00, or_9} + {2'b00, or_14} + {2'b00, or_19} + {2'b00, or_24};

assign sel_decision_0 = {comp_add_0_1 , comp_add_0_1_2_3 , comp_add_0_1_2_3_4};

assign sel_decision_1 = {comp_add_0_1 , comp_add_0_1_2_3 , comp_add_0_1_2_3_4};

assign sel_decision_2 = {comp_add_2_3 , comp_add_0_1_2_3 , comp_add_0_1_2_3_4};

assign sel_decision_3 = {comp_add_2_3 , comp_add_0_1_2_3 , comp_add_0_1_2_3_4};

assign sel_decision_4 = {comp_add_0_1_2_3_4};


	assign comp_add_0_1 = (add_0 >= add_1);
	assign add_0_1 = comp_add_0_1 ? add_0 : add_1;
	assign comp_add_2_3 = (add_2 >= add_3);
	assign add_2_3 = comp_add_2_3 ? add_2 : add_3;
	assign comp_add_0_1_2_3 = (add_0_1 >= add_2_3);
	assign add_0_1_2_3 = comp_add_0_1_2_3 ? add_0_1 : add_2_3;
	assign comp_add_0_1_2_3_4 = (add_0_1_2_3 >= add_4);
	assign add_0_1_2_3_4 = comp_add_0_1_2_3_4 ? add_0_1_2_3 : add_4;
assign reg_decision[0] =  (sel_decision_0 == 3'b111) ? 1'b1 : 1'b0;

assign reg_decision[1] =  (sel_decision_1 == 3'b011) ? 1'b1 : 1'b0;

assign reg_decision[2] =  (sel_decision_2 == 3'b101) ? 1'b1 : 1'b0;

assign reg_decision[3] =  (sel_decision_3 == 3'b001) ? 1'b1 : 1'b0;

assign reg_decision[4] =  (sel_decision_4 == 1'b0) ? 1'b1 : 1'b0;




endmodule
